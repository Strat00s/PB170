/*  Simple 5Khz PWM module
    Start HIGH, stay HIGH until `cnt` = desired_input, reset at after 5000 cycles
*/


module PWM (input clk, input reg[8:0] duty_cycle);
    output out;
    
    initial begin
    
    end

    always @(posedge CLOCK_50) begin


    end

endmodule