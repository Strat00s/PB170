library verilog;
use verilog.vl_types.all;
entity DE2_Default_vlg_vec_tst is
end DE2_Default_vlg_vec_tst;
