library verilog;
use verilog.vl_types.all;
entity knight_rider_vlg_check_tst is
    port(
        clk             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end knight_rider_vlg_check_tst;
