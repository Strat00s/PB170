// system_0.v

// Generated using ACDS version 11.1sp2 259 at 2012.03.31.20:50:59

`timescale 1 ps / 1 ps
module system_0 (
		output wire [9:0]  vga_0_avalon_slave_0_export_VGA_R,        //     vga_0_avalon_slave_0_export.VGA_R
		output wire [9:0]  vga_0_avalon_slave_0_export_VGA_G,        //                                .VGA_G
		output wire [9:0]  vga_0_avalon_slave_0_export_VGA_B,        //                                .VGA_B
		output wire        vga_0_avalon_slave_0_export_VGA_HS,       //                                .VGA_HS
		output wire        vga_0_avalon_slave_0_export_VGA_VS,       //                                .VGA_VS
		output wire        vga_0_avalon_slave_0_export_VGA_SYNC,     //                                .VGA_SYNC
		output wire        vga_0_avalon_slave_0_export_VGA_BLANK,    //                                .VGA_BLANK
		output wire        vga_0_avalon_slave_0_export_VGA_CLK,      //                                .VGA_CLK
		input  wire        vga_0_avalon_slave_0_export_iCLK_25,      //                                .iCLK_25
		input  wire        clk_50,                                   //                   clk_50_clk_in.clk
		inout  wire [3:0]  bidir_port_to_and_from_the_SD_DAT,        //      SD_DAT_external_connection.export
		inout  wire        i2c_sda_external_connection_export,       //     i2c_sda_external_connection.export
		output wire [17:0] out_port_from_the_led_red,                //     led_red_external_connection.export
		input  wire        clk_audio_clk_in_clk,                     //                clk_audio_clk_in.clk
		output wire [6:0]  seg7_display_conduit_end_oSEG0,           //        seg7_display_conduit_end.oSEG0
		output wire [6:0]  seg7_display_conduit_end_oSEG1,           //                                .oSEG1
		output wire [6:0]  seg7_display_conduit_end_oSEG2,           //                                .oSEG2
		output wire [6:0]  seg7_display_conduit_end_oSEG3,           //                                .oSEG3
		output wire [6:0]  seg7_display_conduit_end_oSEG4,           //                                .oSEG4
		output wire [6:0]  seg7_display_conduit_end_oSEG5,           //                                .oSEG5
		output wire [6:0]  seg7_display_conduit_end_oSEG6,           //                                .oSEG6
		output wire [6:0]  seg7_display_conduit_end_oSEG7,           //                                .oSEG7
		output wire [11:0] zs_addr_from_the_sdram_0,                 //                    sdram_0_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram_0,                   //                                .ba
		output wire        zs_cas_n_from_the_sdram_0,                //                                .cas_n
		output wire        zs_cke_from_the_sdram_0,                  //                                .cke
		output wire        zs_cs_n_from_the_sdram_0,                 //                                .cs_n
		inout  wire [15:0] zs_dq_to_and_from_the_sdram_0,            //                                .dq
		output wire [1:0]  zs_dqm_from_the_sdram_0,                  //                                .dqm
		output wire        zs_ras_n_from_the_sdram_0,                //                                .ras_n
		output wire        zs_we_n_from_the_sdram_0,                 //                                .we_n
		input  wire        sd_wp_n_external_connection_export,       //     sd_wp_n_external_connection.export
		inout  wire [7:0]  tri_state_bridge_0_data,                  // tri_state_bridge_0_bridge_0_out.tri_state_bridge_0_data
		output wire        tri_state_bridge_0_readn,                 //                                .tri_state_bridge_0_readn
		output wire        write_n_to_the_cfi_flash_0,               //                                .write_n_to_the_cfi_flash_0
		output wire [21:0] tri_state_bridge_0_address,               //                                .tri_state_bridge_0_address
		output wire        select_n_to_the_cfi_flash_0,              //                                .select_n_to_the_cfi_flash_0
		input  wire        reset_n,                                  //          merged_resets_in_reset.reset_n
		inout  wire        bidir_port_to_and_from_the_SD_CMD,        //      SD_CMD_external_connection.export
		output wire        i2c_scl_external_connection_export,       //     i2c_scl_external_connection.export
		input  wire [3:0]  in_port_to_the_button_pio,                //  button_pio_external_connection.export
		output wire        out_port_from_the_SD_CLK,                 //      SD_CLK_external_connection.export
		inout  wire [15:0] ISP1362_conduit_end_DATA,                 //             ISP1362_conduit_end.DATA
		output wire [1:0]  ISP1362_conduit_end_ADDR,                 //                                .ADDR
		output wire        ISP1362_conduit_end_RD_N,                 //                                .RD_N
		output wire        ISP1362_conduit_end_WR_N,                 //                                .WR_N
		output wire        ISP1362_conduit_end_CS_N,                 //                                .CS_N
		output wire        ISP1362_conduit_end_RST_N,                //                                .RST_N
		input  wire        ISP1362_conduit_end_INT0,                 //                                .INT0
		input  wire        ISP1362_conduit_end_INT1,                 //                                .INT1
		output wire [8:0]  out_port_from_the_led_green,              //   led_green_external_connection.export
		output wire        audio_conduit_end_XCK,                    //               audio_conduit_end.XCK
		input  wire        audio_conduit_end_ADCDAT,                 //                                .ADCDAT
		input  wire        audio_conduit_end_ADCLRC,                 //                                .ADCLRC
		output wire        audio_conduit_end_DACDAT,                 //                                .DACDAT
		input  wire        audio_conduit_end_DACLRC,                 //                                .DACLRC
		input  wire        audio_conduit_end_BCLK,                   //                                .BCLK
		inout  wire [15:0] sram_0_avalon_slave_0_export_DQ,          //    sram_0_avalon_slave_0_export.DQ
		output wire [17:0] sram_0_avalon_slave_0_export_ADDR,        //                                .ADDR
		output wire        sram_0_avalon_slave_0_export_UB_N,        //                                .UB_N
		output wire        sram_0_avalon_slave_0_export_LB_N,        //                                .LB_N
		output wire        sram_0_avalon_slave_0_export_WE_N,        //                                .WE_N
		output wire        sram_0_avalon_slave_0_export_CE_N,        //                                .CE_N
		output wire        sram_0_avalon_slave_0_export_OE_N,        //                                .OE_N
		input  wire        clk,                                      //                      clk_clk_in.clk
		input  wire [17:0] in_port_to_the_switch_pio,                //  switch_pio_external_connection.export
		inout  wire [7:0]  LCD_data_to_and_from_the_lcd_16207_0,     //            lcd_16207_0_external.data
		output wire        LCD_E_from_the_lcd_16207_0,               //                                .E
		output wire        LCD_RS_from_the_lcd_16207_0,              //                                .RS
		output wire        LCD_RW_from_the_lcd_16207_0,              //                                .RW
		input  wire        rxd_to_the_uart_0,                        //      uart_0_external_connection.rxd
		output wire        txd_from_the_uart_0,                      //                                .txd
		input  wire        dm9000a_avalon_slave_0_export_iOSC_50,    //   dm9000a_avalon_slave_0_export.iOSC_50
		inout  wire [15:0] dm9000a_avalon_slave_0_export_ENET_DATA,  //                                .ENET_DATA
		output wire        dm9000a_avalon_slave_0_export_ENET_CMD,   //                                .ENET_CMD
		output wire        dm9000a_avalon_slave_0_export_ENET_RD_N,  //                                .ENET_RD_N
		output wire        dm9000a_avalon_slave_0_export_ENET_WR_N,  //                                .ENET_WR_N
		output wire        dm9000a_avalon_slave_0_export_ENET_CS_N,  //                                .ENET_CS_N
		output wire        dm9000a_avalon_slave_0_export_ENET_RST_N, //                                .ENET_RST_N
		output wire        dm9000a_avalon_slave_0_export_ENET_CLK,   //                                .ENET_CLK
		input  wire        dm9000a_avalon_slave_0_export_ENET_INT    //                                .ENET_INT
	);

	wire   [0:0] tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out;                                     // tri_state_bridge_0_pinSharer_0:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_select_n_to_the_cfi_flash_0
	wire  [21:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out;                                      // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_address -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_address
	wire         tri_state_bridge_0_pinsharer_0_tcm_grant;                                                               // tri_state_bridge_0_bridge_0:grant -> tri_state_bridge_0_pinSharer_0:grant
	wire   [0:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out;                                        // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_readn -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_readn
	wire         tri_state_bridge_0_pinsharer_0_tcm_request;                                                             // tri_state_bridge_0_pinSharer_0:request -> tri_state_bridge_0_bridge_0:request
	wire   [7:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in;                                          // tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_in -> tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_in
	wire         tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen;                                       // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_outen -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_outen
	wire   [0:0] tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out;                                      // tri_state_bridge_0_pinSharer_0:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_write_n_to_the_cfi_flash_0
	wire   [7:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out;                                         // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data
	wire         cfi_flash_0_tcm_chipselect_n_out;                                                                       // cfi_flash_0:tcm_chipselect_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_chipselect_n_out
	wire         cfi_flash_0_tcm_grant;                                                                                  // tri_state_bridge_0_pinSharer_0:tcs0_grant -> cfi_flash_0:tcm_grant
	wire         cfi_flash_0_tcm_data_outen;                                                                             // cfi_flash_0:tcm_data_outen -> tri_state_bridge_0_pinSharer_0:tcs0_data_outen
	wire         cfi_flash_0_tcm_request;                                                                                // cfi_flash_0:tcm_request -> tri_state_bridge_0_pinSharer_0:tcs0_request
	wire   [7:0] cfi_flash_0_tcm_data_out;                                                                               // cfi_flash_0:tcm_data_out -> tri_state_bridge_0_pinSharer_0:tcs0_data_out
	wire         cfi_flash_0_tcm_write_n_out;                                                                            // cfi_flash_0:tcm_write_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_write_n_out
	wire  [21:0] cfi_flash_0_tcm_address_out;                                                                            // cfi_flash_0:tcm_address_out -> tri_state_bridge_0_pinSharer_0:tcs0_address_out
	wire   [7:0] cfi_flash_0_tcm_data_in;                                                                                // tri_state_bridge_0_pinSharer_0:tcs0_data_in -> cfi_flash_0:tcm_data_in
	wire         cfi_flash_0_tcm_read_n_out;                                                                             // cfi_flash_0:tcm_read_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_read_n_out
	wire         cpu_0_instruction_master_waitrequest;                                                                   // cpu_0_instruction_master_translator:av_waitrequest -> cpu_0:i_waitrequest
	wire  [24:0] cpu_0_instruction_master_address;                                                                       // cpu_0:i_address -> cpu_0_instruction_master_translator:av_address
	wire         cpu_0_instruction_master_read;                                                                          // cpu_0:i_read -> cpu_0_instruction_master_translator:av_read
	wire  [31:0] cpu_0_instruction_master_readdata;                                                                      // cpu_0_instruction_master_translator:av_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_readdatavalid;                                                                 // cpu_0_instruction_master_translator:av_readdatavalid -> cpu_0:i_readdatavalid
	wire         cpu_0_data_master_waitrequest;                                                                          // cpu_0_data_master_translator:av_waitrequest -> cpu_0:d_waitrequest
	wire  [31:0] cpu_0_data_master_writedata;                                                                            // cpu_0:d_writedata -> cpu_0_data_master_translator:av_writedata
	wire  [24:0] cpu_0_data_master_address;                                                                              // cpu_0:d_address -> cpu_0_data_master_translator:av_address
	wire         cpu_0_data_master_write;                                                                                // cpu_0:d_write -> cpu_0_data_master_translator:av_write
	wire         cpu_0_data_master_read;                                                                                 // cpu_0:d_read -> cpu_0_data_master_translator:av_read
	wire  [31:0] cpu_0_data_master_readdata;                                                                             // cpu_0_data_master_translator:av_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_debugaccess;                                                                          // cpu_0:jtag_debug_module_debugaccess_to_roms -> cpu_0_data_master_translator:av_debugaccess
	wire   [3:0] cpu_0_data_master_byteenable;                                                                           // cpu_0:d_byteenable -> cpu_0_data_master_translator:av_byteenable
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                       // cpu_0_jtag_debug_module_translator:av_writedata -> cpu_0:jtag_debug_module_writedata
	wire   [8:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                         // cpu_0_jtag_debug_module_translator:av_address -> cpu_0:jtag_debug_module_address
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                      // cpu_0_jtag_debug_module_translator:av_chipselect -> cpu_0:jtag_debug_module_select
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                           // cpu_0_jtag_debug_module_translator:av_write -> cpu_0:jtag_debug_module_write
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                        // cpu_0:jtag_debug_module_readdata -> cpu_0_jtag_debug_module_translator:av_readdata
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                   // cpu_0_jtag_debug_module_translator:av_begintransfer -> cpu_0:jtag_debug_module_begintransfer
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                     // cpu_0_jtag_debug_module_translator:av_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire   [3:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                      // cpu_0_jtag_debug_module_translator:av_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire         sdram_0_s1_translator_avalon_anti_slave_0_waitrequest;                                                  // sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	wire  [15:0] sdram_0_s1_translator_avalon_anti_slave_0_writedata;                                                    // sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	wire  [21:0] sdram_0_s1_translator_avalon_anti_slave_0_address;                                                      // sdram_0_s1_translator:av_address -> sdram_0:az_addr
	wire         sdram_0_s1_translator_avalon_anti_slave_0_chipselect;                                                   // sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	wire         sdram_0_s1_translator_avalon_anti_slave_0_write;                                                        // sdram_0_s1_translator:av_write -> sdram_0:az_wr_n
	wire         sdram_0_s1_translator_avalon_anti_slave_0_read;                                                         // sdram_0_s1_translator:av_read -> sdram_0:az_rd_n
	wire  [15:0] sdram_0_s1_translator_avalon_anti_slave_0_readdata;                                                     // sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	wire         sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid;                                                // sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	wire   [1:0] sdram_0_s1_translator_avalon_anti_slave_0_byteenable;                                                   // sdram_0_s1_translator:av_byteenable -> sdram_0:az_be_n
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata;                             // epcs_controller_epcs_control_port_translator:av_writedata -> epcs_controller:writedata
	wire   [8:0] epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address;                               // epcs_controller_epcs_control_port_translator:av_address -> epcs_controller:address
	wire         epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect;                            // epcs_controller_epcs_control_port_translator:av_chipselect -> epcs_controller:chipselect
	wire         epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write;                                 // epcs_controller_epcs_control_port_translator:av_write -> epcs_controller:write_n
	wire         epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read;                                  // epcs_controller_epcs_control_port_translator:av_read -> epcs_controller:read_n
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata;                              // epcs_controller:readdata -> epcs_controller_epcs_control_port_translator:av_readdata
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest;                                             // cfi_flash_0:uas_waitrequest -> cfi_flash_0_uas_translator:av_waitrequest
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount;                                              // cfi_flash_0_uas_translator:av_burstcount -> cfi_flash_0:uas_burstcount
	wire   [7:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata;                                               // cfi_flash_0_uas_translator:av_writedata -> cfi_flash_0:uas_writedata
	wire  [21:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_address;                                                 // cfi_flash_0_uas_translator:av_address -> cfi_flash_0:uas_address
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_lock;                                                    // cfi_flash_0_uas_translator:av_lock -> cfi_flash_0:uas_lock
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_write;                                                   // cfi_flash_0_uas_translator:av_write -> cfi_flash_0:uas_write
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_read;                                                    // cfi_flash_0_uas_translator:av_read -> cfi_flash_0:uas_read
	wire   [7:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata;                                                // cfi_flash_0:uas_readdata -> cfi_flash_0_uas_translator:av_readdata
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess;                                             // cfi_flash_0_uas_translator:av_debugaccess -> cfi_flash_0:uas_debugaccess
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid;                                           // cfi_flash_0:uas_readdatavalid -> cfi_flash_0_uas_translator:av_readdatavalid
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable;                                              // cfi_flash_0_uas_translator:av_byteenable -> cfi_flash_0:uas_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                               // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                 // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                     // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                      // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                  // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] uart_0_s1_translator_avalon_anti_slave_0_writedata;                                                     // uart_0_s1_translator:av_writedata -> uart_0:writedata
	wire   [2:0] uart_0_s1_translator_avalon_anti_slave_0_address;                                                       // uart_0_s1_translator:av_address -> uart_0:address
	wire         uart_0_s1_translator_avalon_anti_slave_0_chipselect;                                                    // uart_0_s1_translator:av_chipselect -> uart_0:chipselect
	wire         uart_0_s1_translator_avalon_anti_slave_0_write;                                                         // uart_0_s1_translator:av_write -> uart_0:write_n
	wire         uart_0_s1_translator_avalon_anti_slave_0_read;                                                          // uart_0_s1_translator:av_read -> uart_0:read_n
	wire  [15:0] uart_0_s1_translator_avalon_anti_slave_0_readdata;                                                      // uart_0:readdata -> uart_0_s1_translator:av_readdata
	wire         uart_0_s1_translator_avalon_anti_slave_0_begintransfer;                                                 // uart_0_s1_translator:av_begintransfer -> uart_0:begintransfer
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                      // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                        // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire  [15:0] timer_1_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_1_s1_translator:av_writedata -> timer_1:writedata
	wire   [2:0] timer_1_s1_translator_avalon_anti_slave_0_address;                                                      // timer_1_s1_translator:av_address -> timer_1:address
	wire         timer_1_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	wire         timer_1_s1_translator_avalon_anti_slave_0_write;                                                        // timer_1_s1_translator:av_write -> timer_1:write_n
	wire  [15:0] timer_1_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_1:readdata -> timer_1_s1_translator:av_readdata
	wire   [7:0] lcd_control_slave_translator_avalon_anti_slave_0_writedata;                                             // lcd_control_slave_translator:av_writedata -> lcd:writedata
	wire   [1:0] lcd_control_slave_translator_avalon_anti_slave_0_address;                                               // lcd_control_slave_translator:av_address -> lcd:address
	wire         lcd_control_slave_translator_avalon_anti_slave_0_write;                                                 // lcd_control_slave_translator:av_write -> lcd:write
	wire         lcd_control_slave_translator_avalon_anti_slave_0_read;                                                  // lcd_control_slave_translator:av_read -> lcd:read
	wire   [7:0] lcd_control_slave_translator_avalon_anti_slave_0_readdata;                                              // lcd:readdata -> lcd_control_slave_translator:av_readdata
	wire         lcd_control_slave_translator_avalon_anti_slave_0_begintransfer;                                         // lcd_control_slave_translator:av_begintransfer -> lcd:begintransfer
	wire  [31:0] ledr_s1_translator_avalon_anti_slave_0_writedata;                                                       // ledr_s1_translator:av_writedata -> ledr:writedata
	wire   [1:0] ledr_s1_translator_avalon_anti_slave_0_address;                                                         // ledr_s1_translator:av_address -> ledr:address
	wire         ledr_s1_translator_avalon_anti_slave_0_chipselect;                                                      // ledr_s1_translator:av_chipselect -> ledr:chipselect
	wire         ledr_s1_translator_avalon_anti_slave_0_write;                                                           // ledr_s1_translator:av_write -> ledr:write_n
	wire  [31:0] ledr_s1_translator_avalon_anti_slave_0_readdata;                                                        // ledr:readdata -> ledr_s1_translator:av_readdata
	wire  [31:0] ledg_s1_translator_avalon_anti_slave_0_writedata;                                                       // ledg_s1_translator:av_writedata -> ledg:writedata
	wire   [1:0] ledg_s1_translator_avalon_anti_slave_0_address;                                                         // ledg_s1_translator:av_address -> ledg:address
	wire         ledg_s1_translator_avalon_anti_slave_0_chipselect;                                                      // ledg_s1_translator:av_chipselect -> ledg:chipselect
	wire         ledg_s1_translator_avalon_anti_slave_0_write;                                                           // ledg_s1_translator:av_write -> ledg:write_n
	wire  [31:0] ledg_s1_translator_avalon_anti_slave_0_readdata;                                                        // ledg:readdata -> ledg_s1_translator:av_readdata
	wire  [31:0] button_pio_s1_translator_avalon_anti_slave_0_writedata;                                                 // button_pio_s1_translator:av_writedata -> button_pio:writedata
	wire   [1:0] button_pio_s1_translator_avalon_anti_slave_0_address;                                                   // button_pio_s1_translator:av_address -> button_pio:address
	wire         button_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                // button_pio_s1_translator:av_chipselect -> button_pio:chipselect
	wire         button_pio_s1_translator_avalon_anti_slave_0_write;                                                     // button_pio_s1_translator:av_write -> button_pio:write_n
	wire  [31:0] button_pio_s1_translator_avalon_anti_slave_0_readdata;                                                  // button_pio:readdata -> button_pio_s1_translator:av_readdata
	wire   [1:0] switch_pio_s1_translator_avalon_anti_slave_0_address;                                                   // switch_pio_s1_translator:av_address -> switch_pio:address
	wire  [31:0] switch_pio_s1_translator_avalon_anti_slave_0_readdata;                                                  // switch_pio:readdata -> switch_pio_s1_translator:av_readdata
	wire  [31:0] sd_dat_s1_translator_avalon_anti_slave_0_writedata;                                                     // SD_DAT_s1_translator:av_writedata -> SD_DAT:writedata
	wire   [1:0] sd_dat_s1_translator_avalon_anti_slave_0_address;                                                       // SD_DAT_s1_translator:av_address -> SD_DAT:address
	wire         sd_dat_s1_translator_avalon_anti_slave_0_chipselect;                                                    // SD_DAT_s1_translator:av_chipselect -> SD_DAT:chipselect
	wire         sd_dat_s1_translator_avalon_anti_slave_0_write;                                                         // SD_DAT_s1_translator:av_write -> SD_DAT:write_n
	wire  [31:0] sd_dat_s1_translator_avalon_anti_slave_0_readdata;                                                      // SD_DAT:readdata -> SD_DAT_s1_translator:av_readdata
	wire  [31:0] sd_cmd_s1_translator_avalon_anti_slave_0_writedata;                                                     // SD_CMD_s1_translator:av_writedata -> SD_CMD:writedata
	wire   [1:0] sd_cmd_s1_translator_avalon_anti_slave_0_address;                                                       // SD_CMD_s1_translator:av_address -> SD_CMD:address
	wire         sd_cmd_s1_translator_avalon_anti_slave_0_chipselect;                                                    // SD_CMD_s1_translator:av_chipselect -> SD_CMD:chipselect
	wire         sd_cmd_s1_translator_avalon_anti_slave_0_write;                                                         // SD_CMD_s1_translator:av_write -> SD_CMD:write_n
	wire  [31:0] sd_cmd_s1_translator_avalon_anti_slave_0_readdata;                                                      // SD_CMD:readdata -> SD_CMD_s1_translator:av_readdata
	wire  [31:0] sd_clk_s1_translator_avalon_anti_slave_0_writedata;                                                     // SD_CLK_s1_translator:av_writedata -> SD_CLK:writedata
	wire   [1:0] sd_clk_s1_translator_avalon_anti_slave_0_address;                                                       // SD_CLK_s1_translator:av_address -> SD_CLK:address
	wire         sd_clk_s1_translator_avalon_anti_slave_0_chipselect;                                                    // SD_CLK_s1_translator:av_chipselect -> SD_CLK:chipselect
	wire         sd_clk_s1_translator_avalon_anti_slave_0_write;                                                         // SD_CLK_s1_translator:av_write -> SD_CLK:write_n
	wire  [31:0] sd_clk_s1_translator_avalon_anti_slave_0_readdata;                                                      // SD_CLK:readdata -> SD_CLK_s1_translator:av_readdata
	wire  [15:0] isp1362_dc_translator_avalon_anti_slave_0_writedata;                                                    // ISP1362_dc_translator:av_writedata -> ISP1362:avs_dc_writedata_iDATA
	wire         isp1362_dc_translator_avalon_anti_slave_0_address;                                                      // ISP1362_dc_translator:av_address -> ISP1362:avs_dc_address_iADDR
	wire         isp1362_dc_translator_avalon_anti_slave_0_chipselect;                                                   // ISP1362_dc_translator:av_chipselect -> ISP1362:avs_dc_chipselect_n_iCS_N
	wire         isp1362_dc_translator_avalon_anti_slave_0_write;                                                        // ISP1362_dc_translator:av_write -> ISP1362:avs_dc_write_n_iWR_N
	wire         isp1362_dc_translator_avalon_anti_slave_0_read;                                                         // ISP1362_dc_translator:av_read -> ISP1362:avs_dc_read_n_iRD_N
	wire  [15:0] isp1362_dc_translator_avalon_anti_slave_0_readdata;                                                     // ISP1362:avs_dc_readdata_oDATA -> ISP1362_dc_translator:av_readdata
	wire  [15:0] isp1362_hc_translator_avalon_anti_slave_0_writedata;                                                    // ISP1362_hc_translator:av_writedata -> ISP1362:avs_hc_writedata_iDATA
	wire         isp1362_hc_translator_avalon_anti_slave_0_address;                                                      // ISP1362_hc_translator:av_address -> ISP1362:avs_hc_address_iADDR
	wire         isp1362_hc_translator_avalon_anti_slave_0_chipselect;                                                   // ISP1362_hc_translator:av_chipselect -> ISP1362:avs_hc_chipselect_n_iCS_N
	wire         isp1362_hc_translator_avalon_anti_slave_0_write;                                                        // ISP1362_hc_translator:av_write -> ISP1362:avs_hc_write_n_iWR_N
	wire         isp1362_hc_translator_avalon_anti_slave_0_read;                                                         // ISP1362_hc_translator:av_read -> ISP1362:avs_hc_read_n_iRD_N
	wire  [15:0] isp1362_hc_translator_avalon_anti_slave_0_readdata;                                                     // ISP1362:avs_hc_readdata_oDATA -> ISP1362_hc_translator:av_readdata
	wire  [15:0] vga_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                          // VGA_0_avalon_slave_0_translator:av_writedata -> VGA_0:iDATA
	wire  [18:0] vga_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                            // VGA_0_avalon_slave_0_translator:av_address -> VGA_0:iADDR
	wire         vga_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                         // VGA_0_avalon_slave_0_translator:av_chipselect -> VGA_0:iCS
	wire         vga_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                              // VGA_0_avalon_slave_0_translator:av_write -> VGA_0:iWR
	wire         vga_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                               // VGA_0_avalon_slave_0_translator:av_read -> VGA_0:iRD
	wire  [15:0] vga_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                           // VGA_0:oDATA -> VGA_0_avalon_slave_0_translator:av_readdata
	wire  [15:0] dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                        // DM9000A_avalon_slave_0_translator:av_writedata -> DM9000A:iDATA
	wire         dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address;                                          // DM9000A_avalon_slave_0_translator:av_address -> DM9000A:iCMD
	wire         dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                       // DM9000A_avalon_slave_0_translator:av_chipselect -> DM9000A:iCS_N
	wire         dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write;                                            // DM9000A_avalon_slave_0_translator:av_write -> DM9000A:iWR_N
	wire         dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read;                                             // DM9000A_avalon_slave_0_translator:av_read -> DM9000A:iRD_N
	wire  [15:0] dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                         // DM9000A:oDATA -> DM9000A_avalon_slave_0_translator:av_readdata
	wire  [31:0] seg7_avalon_slave_translator_avalon_anti_slave_0_writedata;                                             // seg7_avalon_slave_translator:av_writedata -> seg7:iDIG
	wire         seg7_avalon_slave_translator_avalon_anti_slave_0_write;                                                 // seg7_avalon_slave_translator:av_write -> seg7:iWR
	wire  [15:0] sram_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                         // sram_0_avalon_slave_0_translator:av_writedata -> sram_0:iDATA
	wire  [17:0] sram_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                           // sram_0_avalon_slave_0_translator:av_address -> sram_0:iADDR
	wire         sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                        // sram_0_avalon_slave_0_translator:av_chipselect -> sram_0:iCE_N
	wire         sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                             // sram_0_avalon_slave_0_translator:av_write -> sram_0:iWE_N
	wire         sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                              // sram_0_avalon_slave_0_translator:av_read -> sram_0:iOE_N
	wire  [15:0] sram_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                          // sram_0:oDATA -> sram_0_avalon_slave_0_translator:av_readdata
	wire   [1:0] sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                        // sram_0_avalon_slave_0_translator:av_byteenable -> sram_0:iBE_N
	wire  [31:0] i2c_sda_s1_translator_avalon_anti_slave_0_writedata;                                                    // i2c_sda_s1_translator:av_writedata -> i2c_sda:writedata
	wire   [1:0] i2c_sda_s1_translator_avalon_anti_slave_0_address;                                                      // i2c_sda_s1_translator:av_address -> i2c_sda:address
	wire         i2c_sda_s1_translator_avalon_anti_slave_0_chipselect;                                                   // i2c_sda_s1_translator:av_chipselect -> i2c_sda:chipselect
	wire         i2c_sda_s1_translator_avalon_anti_slave_0_write;                                                        // i2c_sda_s1_translator:av_write -> i2c_sda:write_n
	wire  [31:0] i2c_sda_s1_translator_avalon_anti_slave_0_readdata;                                                     // i2c_sda:readdata -> i2c_sda_s1_translator:av_readdata
	wire  [31:0] i2c_scl_s1_translator_avalon_anti_slave_0_writedata;                                                    // i2c_scl_s1_translator:av_writedata -> i2c_scl:writedata
	wire   [1:0] i2c_scl_s1_translator_avalon_anti_slave_0_address;                                                      // i2c_scl_s1_translator:av_address -> i2c_scl:address
	wire         i2c_scl_s1_translator_avalon_anti_slave_0_chipselect;                                                   // i2c_scl_s1_translator:av_chipselect -> i2c_scl:chipselect
	wire         i2c_scl_s1_translator_avalon_anti_slave_0_write;                                                        // i2c_scl_s1_translator:av_write -> i2c_scl:write_n
	wire  [31:0] i2c_scl_s1_translator_avalon_anti_slave_0_readdata;                                                     // i2c_scl:readdata -> i2c_scl_s1_translator:av_readdata
	wire   [1:0] sd_wp_n_s1_translator_avalon_anti_slave_0_address;                                                      // sd_wp_n_s1_translator:av_address -> sd_wp_n:address
	wire  [31:0] sd_wp_n_s1_translator_avalon_anti_slave_0_readdata;                                                     // sd_wp_n:readdata -> sd_wp_n_s1_translator:av_readdata
	wire  [15:0] audio_avalon_slave_translator_avalon_anti_slave_0_writedata;                                            // audio_avalon_slave_translator:av_writedata -> audio:avs_s1_writedata
	wire   [2:0] audio_avalon_slave_translator_avalon_anti_slave_0_address;                                              // audio_avalon_slave_translator:av_address -> audio:avs_s1_address
	wire         audio_avalon_slave_translator_avalon_anti_slave_0_write;                                                // audio_avalon_slave_translator:av_write -> audio:avs_s1_write
	wire         audio_avalon_slave_translator_avalon_anti_slave_0_read;                                                 // audio_avalon_slave_translator:av_read -> audio:avs_s1_read
	wire  [15:0] audio_avalon_slave_translator_avalon_anti_slave_0_readdata;                                             // audio:avs_s1_readdata -> audio_avalon_slave_translator:av_readdata
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // lcd_control_slave_translator:uav_waitrequest -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_control_slave_translator:uav_burstcount
	wire  [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                               // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_control_slave_translator:uav_writedata
	wire  [24:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                                 // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> lcd_control_slave_translator:uav_address
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                   // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> lcd_control_slave_translator:uav_write
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                    // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_control_slave_translator:uav_lock
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                    // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> lcd_control_slave_translator:uav_read
	wire  [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                // lcd_control_slave_translator:uav_readdata -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // lcd_control_slave_translator:uav_readdatavalid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_control_slave_translator:uav_debugaccess
	wire   [3:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_control_slave_translator:uav_byteenable
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                             // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // ISP1362_hc_translator:uav_waitrequest -> ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] isp1362_hc_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_burstcount -> ISP1362_hc_translator:uav_burstcount
	wire  [31:0] isp1362_hc_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_writedata -> ISP1362_hc_translator:uav_writedata
	wire  [24:0] isp1362_hc_translator_avalon_universal_slave_0_agent_m0_address;                                        // ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_address -> ISP1362_hc_translator:uav_address
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_m0_write;                                          // ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_write -> ISP1362_hc_translator:uav_write
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_m0_lock;                                           // ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_lock -> ISP1362_hc_translator:uav_lock
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_m0_read;                                           // ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_read -> ISP1362_hc_translator:uav_read
	wire  [31:0] isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // ISP1362_hc_translator:uav_readdata -> ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // ISP1362_hc_translator:uav_readdatavalid -> ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ISP1362_hc_translator:uav_debugaccess
	wire   [3:0] isp1362_hc_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_byteenable -> ISP1362_hc_translator:uav_byteenable
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_valid -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_data -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // sd_wp_n_s1_translator:uav_waitrequest -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sd_wp_n_s1_translator:uav_burstcount
	wire  [31:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sd_wp_n_s1_translator:uav_writedata
	wire  [24:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_address -> sd_wp_n_s1_translator:uav_address
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_write -> sd_wp_n_s1_translator:uav_write
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sd_wp_n_s1_translator:uav_lock
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_read -> sd_wp_n_s1_translator:uav_read
	wire  [31:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // sd_wp_n_s1_translator:uav_readdata -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // sd_wp_n_s1_translator:uav_readdatavalid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sd_wp_n_s1_translator:uav_debugaccess
	wire   [3:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sd_wp_n_s1_translator:uav_byteenable
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [24:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // switch_pio_s1_translator:uav_waitrequest -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch_pio_s1_translator:uav_burstcount
	wire  [31:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch_pio_s1_translator:uav_writedata
	wire  [24:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch_pio_s1_translator:uav_address
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch_pio_s1_translator:uav_write
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch_pio_s1_translator:uav_lock
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch_pio_s1_translator:uav_read
	wire  [31:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // switch_pio_s1_translator:uav_readdata -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // switch_pio_s1_translator:uav_readdatavalid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch_pio_s1_translator:uav_debugaccess
	wire   [3:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch_pio_s1_translator:uav_byteenable
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // ledg_s1_translator:uav_waitrequest -> ledg_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // ledg_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ledg_s1_translator:uav_burstcount
	wire  [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // ledg_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ledg_s1_translator:uav_writedata
	wire  [24:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // ledg_s1_translator_avalon_universal_slave_0_agent:m0_address -> ledg_s1_translator:uav_address
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // ledg_s1_translator_avalon_universal_slave_0_agent:m0_write -> ledg_s1_translator:uav_write
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // ledg_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ledg_s1_translator:uav_lock
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // ledg_s1_translator_avalon_universal_slave_0_agent:m0_read -> ledg_s1_translator:uav_read
	wire  [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // ledg_s1_translator:uav_readdata -> ledg_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // ledg_s1_translator:uav_readdatavalid -> ledg_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // ledg_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ledg_s1_translator:uav_debugaccess
	wire   [3:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // ledg_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ledg_s1_translator:uav_byteenable
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // i2c_sda_s1_translator:uav_waitrequest -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> i2c_sda_s1_translator:uav_burstcount
	wire  [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> i2c_sda_s1_translator:uav_writedata
	wire  [24:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_address -> i2c_sda_s1_translator:uav_address
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_write -> i2c_sda_s1_translator:uav_write
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_lock -> i2c_sda_s1_translator:uav_lock
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_read -> i2c_sda_s1_translator:uav_read
	wire  [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // i2c_sda_s1_translator:uav_readdata -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // i2c_sda_s1_translator:uav_readdatavalid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> i2c_sda_s1_translator:uav_debugaccess
	wire   [3:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> i2c_sda_s1_translator:uav_byteenable
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // button_pio_s1_translator:uav_waitrequest -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_pio_s1_translator:uav_burstcount
	wire  [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_pio_s1_translator:uav_writedata
	wire  [24:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_pio_s1_translator:uav_address
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_pio_s1_translator:uav_write
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_pio_s1_translator:uav_lock
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_pio_s1_translator:uav_read
	wire  [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // button_pio_s1_translator:uav_readdata -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // button_pio_s1_translator:uav_readdatavalid -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_pio_s1_translator:uav_debugaccess
	wire   [3:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_pio_s1_translator:uav_byteenable
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // cpu_0_jtag_debug_module_translator:uav_waitrequest -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_0_jtag_debug_module_translator:uav_writedata
	wire  [24:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                           // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_0_jtag_debug_module_translator:uav_address
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_0_jtag_debug_module_translator:uav_write
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                              // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_0_jtag_debug_module_translator:uav_lock
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                              // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_0_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                          // cpu_0_jtag_debug_module_translator:uav_readdata -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // cpu_0_jtag_debug_module_translator:uav_readdatavalid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_0_jtag_debug_module_translator:uav_byteenable
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // ledr_s1_translator:uav_waitrequest -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // ledr_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ledr_s1_translator:uav_burstcount
	wire  [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // ledr_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ledr_s1_translator:uav_writedata
	wire  [24:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // ledr_s1_translator_avalon_universal_slave_0_agent:m0_address -> ledr_s1_translator:uav_address
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // ledr_s1_translator_avalon_universal_slave_0_agent:m0_write -> ledr_s1_translator:uav_write
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // ledr_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ledr_s1_translator:uav_lock
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // ledr_s1_translator_avalon_universal_slave_0_agent:m0_read -> ledr_s1_translator:uav_read
	wire  [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // ledr_s1_translator:uav_readdata -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // ledr_s1_translator:uav_readdatavalid -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // ledr_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ledr_s1_translator:uav_debugaccess
	wire   [3:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // ledr_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ledr_s1_translator:uav_byteenable
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // seg7_avalon_slave_translator:uav_waitrequest -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> seg7_avalon_slave_translator:uav_burstcount
	wire  [31:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                               // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> seg7_avalon_slave_translator:uav_writedata
	wire  [24:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                                 // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> seg7_avalon_slave_translator:uav_address
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                                   // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> seg7_avalon_slave_translator:uav_write
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                    // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> seg7_avalon_slave_translator:uav_lock
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                                    // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> seg7_avalon_slave_translator:uav_read
	wire  [31:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                // seg7_avalon_slave_translator:uav_readdata -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // seg7_avalon_slave_translator:uav_readdatavalid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seg7_avalon_slave_translator:uav_debugaccess
	wire   [3:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> seg7_avalon_slave_translator:uav_byteenable
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                             // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // cfi_flash_0_uas_translator:uav_waitrequest -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> cfi_flash_0_uas_translator:uav_burstcount
	wire   [7:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> cfi_flash_0_uas_translator:uav_writedata
	wire  [24:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address;                                   // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_address -> cfi_flash_0_uas_translator:uav_address
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write;                                     // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_write -> cfi_flash_0_uas_translator:uav_write
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_lock -> cfi_flash_0_uas_translator:uav_lock
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read;                                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_read -> cfi_flash_0_uas_translator:uav_read
	wire   [7:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // cfi_flash_0_uas_translator:uav_readdata -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // cfi_flash_0_uas_translator:uav_readdatavalid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cfi_flash_0_uas_translator:uav_debugaccess
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> cfi_flash_0_uas_translator:uav_byteenable
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [57:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                               // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [57:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	wire  [24:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	wire   [3:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // SD_CMD_s1_translator:uav_waitrequest -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_CMD_s1_translator:uav_burstcount
	wire  [31:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_CMD_s1_translator:uav_writedata
	wire  [24:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_address -> SD_CMD_s1_translator:uav_address
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_write -> SD_CMD_s1_translator:uav_write
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SD_CMD_s1_translator:uav_lock
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_read -> SD_CMD_s1_translator:uav_read
	wire  [31:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // SD_CMD_s1_translator:uav_readdata -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // SD_CMD_s1_translator:uav_readdatavalid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_CMD_s1_translator:uav_debugaccess
	wire   [3:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_CMD_s1_translator:uav_byteenable
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // uart_0_s1_translator:uav_waitrequest -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_0_s1_translator:uav_burstcount
	wire  [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_0_s1_translator:uav_writedata
	wire  [24:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_0_s1_translator:uav_address
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_0_s1_translator:uav_write
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_0_s1_translator:uav_lock
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_0_s1_translator:uav_read
	wire  [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // uart_0_s1_translator:uav_readdata -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // uart_0_s1_translator:uav_readdatavalid -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_0_s1_translator:uav_debugaccess
	wire   [3:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_0_s1_translator:uav_byteenable
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // DM9000A_avalon_slave_0_translator:uav_waitrequest -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> DM9000A_avalon_slave_0_translator:uav_burstcount
	wire  [31:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                          // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> DM9000A_avalon_slave_0_translator:uav_writedata
	wire  [24:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                            // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> DM9000A_avalon_slave_0_translator:uav_address
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                              // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> DM9000A_avalon_slave_0_translator:uav_write
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                               // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> DM9000A_avalon_slave_0_translator:uav_lock
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                               // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> DM9000A_avalon_slave_0_translator:uav_read
	wire  [31:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                           // DM9000A_avalon_slave_0_translator:uav_readdata -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // DM9000A_avalon_slave_0_translator:uav_readdatavalid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DM9000A_avalon_slave_0_translator:uav_debugaccess
	wire   [3:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> DM9000A_avalon_slave_0_translator:uav_byteenable
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                        // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // ISP1362_dc_translator:uav_waitrequest -> ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] isp1362_dc_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_burstcount -> ISP1362_dc_translator:uav_burstcount
	wire  [31:0] isp1362_dc_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_writedata -> ISP1362_dc_translator:uav_writedata
	wire  [24:0] isp1362_dc_translator_avalon_universal_slave_0_agent_m0_address;                                        // ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_address -> ISP1362_dc_translator:uav_address
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_m0_write;                                          // ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_write -> ISP1362_dc_translator:uav_write
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_m0_lock;                                           // ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_lock -> ISP1362_dc_translator:uav_lock
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_m0_read;                                           // ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_read -> ISP1362_dc_translator:uav_read
	wire  [31:0] isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // ISP1362_dc_translator:uav_readdata -> ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // ISP1362_dc_translator:uav_readdatavalid -> ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ISP1362_dc_translator:uav_debugaccess
	wire   [3:0] isp1362_dc_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_byteenable -> ISP1362_dc_translator:uav_byteenable
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_valid -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_data -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // VGA_0_avalon_slave_0_translator:uav_waitrequest -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_0_avalon_slave_0_translator:uav_burstcount
	wire  [31:0] vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                            // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_0_avalon_slave_0_translator:uav_writedata
	wire  [24:0] vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                              // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> VGA_0_avalon_slave_0_translator:uav_address
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> VGA_0_avalon_slave_0_translator:uav_write
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                 // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_0_avalon_slave_0_translator:uav_lock
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                 // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> VGA_0_avalon_slave_0_translator:uav_read
	wire  [31:0] vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                             // VGA_0_avalon_slave_0_translator:uav_readdata -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // VGA_0_avalon_slave_0_translator:uav_readdatavalid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_0_avalon_slave_0_translator:uav_debugaccess
	wire   [3:0] vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_0_avalon_slave_0_translator:uav_byteenable
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                          // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // audio_avalon_slave_translator:uav_waitrequest -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_avalon_slave_translator:uav_burstcount
	wire  [31:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                              // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_avalon_slave_translator:uav_writedata
	wire  [24:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                                // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> audio_avalon_slave_translator:uav_address
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                                  // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> audio_avalon_slave_translator:uav_write
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                   // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> audio_avalon_slave_translator:uav_lock
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                                   // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> audio_avalon_slave_translator:uav_read
	wire  [31:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                               // audio_avalon_slave_translator:uav_readdata -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // audio_avalon_slave_translator:uav_readdatavalid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_avalon_slave_translator:uav_debugaccess
	wire   [3:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // audio_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_avalon_slave_translator:uav_byteenable
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                            // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [31:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                      // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                       // audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                      // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // SD_CLK_s1_translator:uav_waitrequest -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_CLK_s1_translator:uav_burstcount
	wire  [31:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_CLK_s1_translator:uav_writedata
	wire  [24:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_address -> SD_CLK_s1_translator:uav_address
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_write -> SD_CLK_s1_translator:uav_write
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SD_CLK_s1_translator:uav_lock
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_read -> SD_CLK_s1_translator:uav_read
	wire  [31:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // SD_CLK_s1_translator:uav_readdata -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // SD_CLK_s1_translator:uav_readdatavalid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_CLK_s1_translator:uav_debugaccess
	wire   [3:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_CLK_s1_translator:uav_byteenable
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // epcs_controller_epcs_control_port_translator:uav_waitrequest -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;              // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> epcs_controller_epcs_control_port_translator:uav_burstcount
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;               // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> epcs_controller_epcs_control_port_translator:uav_writedata
	wire  [24:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address;                 // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_address -> epcs_controller_epcs_control_port_translator:uav_address
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write;                   // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_write -> epcs_controller_epcs_control_port_translator:uav_write
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> epcs_controller_epcs_control_port_translator:uav_lock
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read;                    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_read -> epcs_controller_epcs_control_port_translator:uav_read
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                // epcs_controller_epcs_control_port_translator:uav_readdata -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // epcs_controller_epcs_control_port_translator:uav_readdatavalid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epcs_controller_epcs_control_port_translator:uav_debugaccess
	wire   [3:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;              // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> epcs_controller_epcs_control_port_translator:uav_byteenable
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;            // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;             // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;            // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_0_data_master_translator_avalon_universal_master_0_waitrequest;                                     // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_0_data_master_translator_avalon_universal_master_0_burstcount;                                      // cpu_0_data_master_translator:uav_burstcount -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_0_data_master_translator_avalon_universal_master_0_writedata;                                       // cpu_0_data_master_translator:uav_writedata -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] cpu_0_data_master_translator_avalon_universal_master_0_address;                                         // cpu_0_data_master_translator:uav_address -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_0_data_master_translator_avalon_universal_master_0_lock;                                            // cpu_0_data_master_translator:uav_lock -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_0_data_master_translator_avalon_universal_master_0_write;                                           // cpu_0_data_master_translator:uav_write -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_0_data_master_translator_avalon_universal_master_0_read;                                            // cpu_0_data_master_translator:uav_read -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_0_data_master_translator_avalon_universal_master_0_readdata;                                        // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_data_master_translator:uav_readdata
	wire         cpu_0_data_master_translator_avalon_universal_master_0_debugaccess;                                     // cpu_0_data_master_translator:uav_debugaccess -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_0_data_master_translator_avalon_universal_master_0_byteenable;                                      // cpu_0_data_master_translator:uav_byteenable -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                   // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_data_master_translator:uav_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [24:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // SD_DAT_s1_translator:uav_waitrequest -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_DAT_s1_translator:uav_burstcount
	wire  [31:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_DAT_s1_translator:uav_writedata
	wire  [24:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_address -> SD_DAT_s1_translator:uav_address
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_write -> SD_DAT_s1_translator:uav_write
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SD_DAT_s1_translator:uav_lock
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_read -> SD_DAT_s1_translator:uav_read
	wire  [31:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // SD_DAT_s1_translator:uav_readdata -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // SD_DAT_s1_translator:uav_readdatavalid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_DAT_s1_translator:uav_debugaccess
	wire   [3:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_DAT_s1_translator:uav_byteenable
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                              // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount;                               // cpu_0_instruction_master_translator:uav_burstcount -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_writedata;                                // cpu_0_instruction_master_translator:uav_writedata -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] cpu_0_instruction_master_translator_avalon_universal_master_0_address;                                  // cpu_0_instruction_master_translator:uav_address -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_lock;                                     // cpu_0_instruction_master_translator:uav_lock -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_write;                                    // cpu_0_instruction_master_translator:uav_write -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_read;                                     // cpu_0_instruction_master_translator:uav_read -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_readdata;                                 // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_instruction_master_translator:uav_readdata
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                              // cpu_0_instruction_master_translator:uav_debugaccess -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable;                               // cpu_0_instruction_master_translator:uav_byteenable -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                            // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_instruction_master_translator:uav_readdatavalid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	wire  [24:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	wire   [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // i2c_scl_s1_translator:uav_waitrequest -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> i2c_scl_s1_translator:uav_burstcount
	wire  [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> i2c_scl_s1_translator:uav_writedata
	wire  [24:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_address -> i2c_scl_s1_translator:uav_address
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_write -> i2c_scl_s1_translator:uav_write
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> i2c_scl_s1_translator:uav_lock
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_read -> i2c_scl_s1_translator:uav_read
	wire  [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // i2c_scl_s1_translator:uav_readdata -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // i2c_scl_s1_translator:uav_readdatavalid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> i2c_scl_s1_translator:uav_debugaccess
	wire   [3:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> i2c_scl_s1_translator:uav_byteenable
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // sram_0_avalon_slave_0_translator:uav_waitrequest -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_0_avalon_slave_0_translator:uav_burstcount
	wire  [15:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                           // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_0_avalon_slave_0_translator:uav_writedata
	wire  [24:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                             // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> sram_0_avalon_slave_0_translator:uav_address
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                               // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> sram_0_avalon_slave_0_translator:uav_write
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> sram_0_avalon_slave_0_translator:uav_lock
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> sram_0_avalon_slave_0_translator:uav_read
	wire  [15:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                            // sram_0_avalon_slave_0_translator:uav_readdata -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // sram_0_avalon_slave_0_translator:uav_readdatavalid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_0_avalon_slave_0_translator:uav_debugaccess
	wire   [1:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_0_avalon_slave_0_translator:uav_byteenable
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                         // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                     // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                           // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                   // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [83:0] cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                            // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                           // addr_router:sink_ready -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                  // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [83:0] cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                   // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router_001:sink_ready -> cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [83:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                              // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router:sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [65:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_001:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                   // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [83:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data;                    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_002:sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                     // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [56:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data;                                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_003:sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [83:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_004:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [83:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_005:sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [83:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_006:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [83:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_007:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                   // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [83:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                    // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_008:sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // ledr_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // ledr_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // ledr_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [83:0] ledr_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // ledr_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_009:sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // ledg_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // ledg_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // ledg_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [83:0] ledg_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // ledg_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_010:sink_ready -> ledg_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [83:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_011:sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [83:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_012:sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [83:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_013:sink_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [83:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_014:sink_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [83:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_015:sink_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rp_valid;                                          // ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [83:0] isp1362_dc_translator_avalon_universal_slave_0_agent_rp_data;                                           // ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire         isp1362_dc_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_016:sink_ready -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_ready
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rp_valid;                                          // ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [83:0] isp1362_hc_translator_avalon_universal_slave_0_agent_rp_data;                                           // ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire         isp1362_hc_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_017:sink_ready -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_ready
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [83:0] vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                 // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire         vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_018:sink_ready -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                              // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [83:0] dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                               // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire         dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_019:sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                   // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [83:0] seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                                    // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire         seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_020:sink_ready -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                               // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [65:0] sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire         sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_021:sink_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [83:0] i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire         i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_022:sink_ready -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire  [83:0] i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire         i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_023:sink_ready -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire  [83:0] sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire         sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_024:sink_ready -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                  // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire  [83:0] audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                                   // audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire         audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_025:sink_ready -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                            // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                                  // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                          // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [83:0] addr_router_src_data;                                                                                   // addr_router:src_data -> limiter:cmd_sink_data
	wire  [25:0] addr_router_src_channel;                                                                                // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                                  // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                            // limiter:rsp_src_endofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                                  // limiter:rsp_src_valid -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                          // limiter:rsp_src_startofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [83:0] limiter_rsp_src_data;                                                                                   // limiter:rsp_src_data -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [25:0] limiter_rsp_src_channel;                                                                                // limiter:rsp_src_channel -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                                  // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         burst_adapter_source0_endofpacket;                                                                      // burst_adapter:source0_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                            // burst_adapter:source0_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                                    // burst_adapter:source0_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [56:0] burst_adapter_source0_data;                                                                             // burst_adapter:source0_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                            // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire  [25:0] burst_adapter_source0_channel;                                                                          // burst_adapter:source0_channel -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_001_source0_endofpacket;                                                                  // burst_adapter_001:source0_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_001_source0_valid;                                                                        // burst_adapter_001:source0_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_001_source0_startofpacket;                                                                // burst_adapter_001:source0_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_001_source0_data;                                                                         // burst_adapter_001:source0_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_001_source0_ready;                                                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire  [25:0] burst_adapter_001_source0_channel;                                                                      // burst_adapter_001:source0_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_002_source0_endofpacket;                                                                  // burst_adapter_002:source0_endofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_002_source0_valid;                                                                        // burst_adapter_002:source0_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_002_source0_startofpacket;                                                                // burst_adapter_002:source0_startofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_002_source0_data;                                                                         // burst_adapter_002:source0_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_002_source0_ready;                                                                        // sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire  [25:0] burst_adapter_002_source0_channel;                                                                      // burst_adapter_002:source0_channel -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                         // rst_controller:reset_out -> [SD_CLK:reset_n, SD_CLK_s1_translator:reset, SD_CLK_s1_translator_avalon_universal_slave_0_agent:reset, SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_CMD:reset_n, SD_CMD_s1_translator:reset, SD_CMD_s1_translator_avalon_universal_slave_0_agent:reset, SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_DAT:reset_n, SD_DAT_s1_translator:reset, SD_DAT_s1_translator_avalon_universal_slave_0_agent:reset, SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, button_pio:reset_n, button_pio_s1_translator:reset, button_pio_s1_translator_avalon_universal_slave_0_agent:reset, button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cfi_flash_0:reset_reset, cfi_flash_0_uas_translator:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cpu_0:reset_n, cpu_0_data_master_translator:reset, cpu_0_data_master_translator_avalon_universal_master_0_agent:reset, cpu_0_instruction_master_translator:reset, cpu_0_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_0_jtag_debug_module_translator:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:out_reset, epcs_controller:reset_n, epcs_controller_epcs_control_port_translator:reset, epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:reset, epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd:reset_n, lcd_control_slave_translator:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ledg:reset_n, ledg_s1_translator:reset, ledg_s1_translator_avalon_universal_slave_0_agent:reset, ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ledr:reset_n, ledr_s1_translator:reset, ledr_s1_translator_avalon_universal_slave_0_agent:reset, ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram_0:reset_n, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch_pio:reset_n, switch_pio_s1_translator:reset, switch_pio_s1_translator_avalon_universal_slave_0_agent:reset, switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1:reset_n, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tri_state_bridge_0_bridge_0:reset, tri_state_bridge_0_pinSharer_0:reset_reset, uart_0:reset_n, uart_0_s1_translator:reset, uart_0_s1_translator_avalon_universal_slave_0_agent:reset, uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire         cpu_0_jtag_debug_module_reset_reset;                                                                    // cpu_0:jtag_debug_module_resetrequest -> rst_controller:reset_in2
	wire         rst_controller_001_reset_out_reset;                                                                     // rst_controller_001:reset_out -> [DM9000A:iRST_N, DM9000A_avalon_slave_0_translator:reset, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ISP1362:avs_dc_reset_n_iRST_N, ISP1362:avs_hc_reset_n_iRST_N, ISP1362_dc_translator:reset, ISP1362_dc_translator_avalon_universal_slave_0_agent:reset, ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ISP1362_hc_translator:reset, ISP1362_hc_translator_avalon_universal_slave_0_agent:reset, ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_0:iRST_N, VGA_0_avalon_slave_0_translator:reset, VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter_002:reset, i2c_scl:reset_n, i2c_scl_s1_translator:reset, i2c_scl_s1_translator_avalon_universal_slave_0_agent:reset, i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, i2c_sda:reset_n, i2c_sda_s1_translator:reset, i2c_sda_s1_translator_avalon_universal_slave_0_agent:reset, i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, sd_wp_n:reset_n, sd_wp_n_s1_translator:reset, sd_wp_n_s1_translator_avalon_universal_slave_0_agent:reset, sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, seg7:iRST_N, seg7_avalon_slave_translator:reset, seg7_avalon_slave_translator_avalon_universal_slave_0_agent:reset, seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sram_0:iRST_N, sram_0_avalon_slave_0_translator:reset, sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter_004:reset, width_adapter_005:reset]
	wire         rst_controller_002_reset_out_reset;                                                                     // rst_controller_002:reset_out -> [audio:avs_s1_reset, audio_avalon_slave_translator:reset, audio_avalon_slave_translator_avalon_universal_slave_0_agent:reset, audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_001:in_reset, id_router_025:reset, rsp_xbar_demux_025:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                        // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                              // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                      // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src0_data;                                                                               // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [25:0] cmd_xbar_demux_src0_channel;                                                                            // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                              // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                        // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                              // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                      // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src1_data;                                                                               // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [25:0] cmd_xbar_demux_src1_channel;                                                                            // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                              // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                        // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                              // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                      // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src2_data;                                                                               // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [25:0] cmd_xbar_demux_src2_channel;                                                                            // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                              // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                        // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                              // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                      // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src3_data;                                                                               // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire  [25:0] cmd_xbar_demux_src3_channel;                                                                            // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                              // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                    // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                          // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                                  // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src0_data;                                                                           // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [25:0] cmd_xbar_demux_001_src0_channel;                                                                        // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                          // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                    // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                          // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                                  // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src1_data;                                                                           // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [25:0] cmd_xbar_demux_001_src1_channel;                                                                        // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                          // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                    // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                          // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                                  // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src2_data;                                                                           // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [25:0] cmd_xbar_demux_001_src2_channel;                                                                        // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                          // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                    // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                          // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                                  // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src3_data;                                                                           // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire  [25:0] cmd_xbar_demux_001_src3_channel;                                                                        // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                          // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                    // cmd_xbar_demux_001:src4_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                          // cmd_xbar_demux_001:src4_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                                  // cmd_xbar_demux_001:src4_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src4_data;                                                                           // cmd_xbar_demux_001:src4_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src4_channel;                                                                        // cmd_xbar_demux_001:src4_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                    // cmd_xbar_demux_001:src5_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                          // cmd_xbar_demux_001:src5_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                                  // cmd_xbar_demux_001:src5_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src5_data;                                                                           // cmd_xbar_demux_001:src5_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src5_channel;                                                                        // cmd_xbar_demux_001:src5_channel -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                    // cmd_xbar_demux_001:src6_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                          // cmd_xbar_demux_001:src6_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                                  // cmd_xbar_demux_001:src6_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src6_data;                                                                           // cmd_xbar_demux_001:src6_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src6_channel;                                                                        // cmd_xbar_demux_001:src6_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                    // cmd_xbar_demux_001:src7_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                          // cmd_xbar_demux_001:src7_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                                  // cmd_xbar_demux_001:src7_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src7_data;                                                                           // cmd_xbar_demux_001:src7_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src7_channel;                                                                        // cmd_xbar_demux_001:src7_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                    // cmd_xbar_demux_001:src8_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                          // cmd_xbar_demux_001:src8_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                                  // cmd_xbar_demux_001:src8_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src8_data;                                                                           // cmd_xbar_demux_001:src8_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src8_channel;                                                                        // cmd_xbar_demux_001:src8_channel -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                                    // cmd_xbar_demux_001:src9_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                          // cmd_xbar_demux_001:src9_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                                  // cmd_xbar_demux_001:src9_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src9_data;                                                                           // cmd_xbar_demux_001:src9_data -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src9_channel;                                                                        // cmd_xbar_demux_001:src9_channel -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                                   // cmd_xbar_demux_001:src10_endofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                         // cmd_xbar_demux_001:src10_valid -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                                 // cmd_xbar_demux_001:src10_startofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src10_data;                                                                          // cmd_xbar_demux_001:src10_data -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src10_channel;                                                                       // cmd_xbar_demux_001:src10_channel -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                                   // cmd_xbar_demux_001:src11_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                         // cmd_xbar_demux_001:src11_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                                 // cmd_xbar_demux_001:src11_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src11_data;                                                                          // cmd_xbar_demux_001:src11_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src11_channel;                                                                       // cmd_xbar_demux_001:src11_channel -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src12_endofpacket;                                                                   // cmd_xbar_demux_001:src12_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src12_valid;                                                                         // cmd_xbar_demux_001:src12_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src12_startofpacket;                                                                 // cmd_xbar_demux_001:src12_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src12_data;                                                                          // cmd_xbar_demux_001:src12_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src12_channel;                                                                       // cmd_xbar_demux_001:src12_channel -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src13_endofpacket;                                                                   // cmd_xbar_demux_001:src13_endofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src13_valid;                                                                         // cmd_xbar_demux_001:src13_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src13_startofpacket;                                                                 // cmd_xbar_demux_001:src13_startofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src13_data;                                                                          // cmd_xbar_demux_001:src13_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src13_channel;                                                                       // cmd_xbar_demux_001:src13_channel -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src14_endofpacket;                                                                   // cmd_xbar_demux_001:src14_endofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src14_valid;                                                                         // cmd_xbar_demux_001:src14_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src14_startofpacket;                                                                 // cmd_xbar_demux_001:src14_startofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src14_data;                                                                          // cmd_xbar_demux_001:src14_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src14_channel;                                                                       // cmd_xbar_demux_001:src14_channel -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src15_endofpacket;                                                                   // cmd_xbar_demux_001:src15_endofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src15_valid;                                                                         // cmd_xbar_demux_001:src15_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src15_startofpacket;                                                                 // cmd_xbar_demux_001:src15_startofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src15_data;                                                                          // cmd_xbar_demux_001:src15_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src15_channel;                                                                       // cmd_xbar_demux_001:src15_channel -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src16_endofpacket;                                                                   // cmd_xbar_demux_001:src16_endofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src16_valid;                                                                         // cmd_xbar_demux_001:src16_valid -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src16_startofpacket;                                                                 // cmd_xbar_demux_001:src16_startofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src16_data;                                                                          // cmd_xbar_demux_001:src16_data -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src16_channel;                                                                       // cmd_xbar_demux_001:src16_channel -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src17_endofpacket;                                                                   // cmd_xbar_demux_001:src17_endofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src17_valid;                                                                         // cmd_xbar_demux_001:src17_valid -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src17_startofpacket;                                                                 // cmd_xbar_demux_001:src17_startofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src17_data;                                                                          // cmd_xbar_demux_001:src17_data -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src17_channel;                                                                       // cmd_xbar_demux_001:src17_channel -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src18_endofpacket;                                                                   // cmd_xbar_demux_001:src18_endofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src18_valid;                                                                         // cmd_xbar_demux_001:src18_valid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src18_startofpacket;                                                                 // cmd_xbar_demux_001:src18_startofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src18_data;                                                                          // cmd_xbar_demux_001:src18_data -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src18_channel;                                                                       // cmd_xbar_demux_001:src18_channel -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src19_endofpacket;                                                                   // cmd_xbar_demux_001:src19_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src19_valid;                                                                         // cmd_xbar_demux_001:src19_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src19_startofpacket;                                                                 // cmd_xbar_demux_001:src19_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src19_data;                                                                          // cmd_xbar_demux_001:src19_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src19_channel;                                                                       // cmd_xbar_demux_001:src19_channel -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src20_endofpacket;                                                                   // cmd_xbar_demux_001:src20_endofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src20_valid;                                                                         // cmd_xbar_demux_001:src20_valid -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src20_startofpacket;                                                                 // cmd_xbar_demux_001:src20_startofpacket -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src20_data;                                                                          // cmd_xbar_demux_001:src20_data -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src20_channel;                                                                       // cmd_xbar_demux_001:src20_channel -> seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src21_endofpacket;                                                                   // cmd_xbar_demux_001:src21_endofpacket -> width_adapter_004:in_endofpacket
	wire         cmd_xbar_demux_001_src21_valid;                                                                         // cmd_xbar_demux_001:src21_valid -> width_adapter_004:in_valid
	wire         cmd_xbar_demux_001_src21_startofpacket;                                                                 // cmd_xbar_demux_001:src21_startofpacket -> width_adapter_004:in_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src21_data;                                                                          // cmd_xbar_demux_001:src21_data -> width_adapter_004:in_data
	wire  [25:0] cmd_xbar_demux_001_src21_channel;                                                                       // cmd_xbar_demux_001:src21_channel -> width_adapter_004:in_channel
	wire         cmd_xbar_demux_001_src22_endofpacket;                                                                   // cmd_xbar_demux_001:src22_endofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src22_valid;                                                                         // cmd_xbar_demux_001:src22_valid -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src22_startofpacket;                                                                 // cmd_xbar_demux_001:src22_startofpacket -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src22_data;                                                                          // cmd_xbar_demux_001:src22_data -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src22_channel;                                                                       // cmd_xbar_demux_001:src22_channel -> i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src23_endofpacket;                                                                   // cmd_xbar_demux_001:src23_endofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src23_valid;                                                                         // cmd_xbar_demux_001:src23_valid -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src23_startofpacket;                                                                 // cmd_xbar_demux_001:src23_startofpacket -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src23_data;                                                                          // cmd_xbar_demux_001:src23_data -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src23_channel;                                                                       // cmd_xbar_demux_001:src23_channel -> i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src24_endofpacket;                                                                   // cmd_xbar_demux_001:src24_endofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src24_valid;                                                                         // cmd_xbar_demux_001:src24_valid -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src24_startofpacket;                                                                 // cmd_xbar_demux_001:src24_startofpacket -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src24_data;                                                                          // cmd_xbar_demux_001:src24_data -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_demux_001_src24_channel;                                                                       // cmd_xbar_demux_001:src24_channel -> sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                        // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                              // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                      // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [83:0] rsp_xbar_demux_src0_data;                                                                               // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [25:0] rsp_xbar_demux_src0_channel;                                                                            // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                              // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                        // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                              // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                      // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [83:0] rsp_xbar_demux_src1_data;                                                                               // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [25:0] rsp_xbar_demux_src1_channel;                                                                            // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                              // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                    // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                          // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                                  // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [83:0] rsp_xbar_demux_001_src0_data;                                                                           // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [25:0] rsp_xbar_demux_001_src0_channel;                                                                        // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                          // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                    // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                          // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                                  // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [83:0] rsp_xbar_demux_001_src1_data;                                                                           // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [25:0] rsp_xbar_demux_001_src1_channel;                                                                        // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                          // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                    // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                          // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                                  // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [83:0] rsp_xbar_demux_002_src0_data;                                                                           // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [25:0] rsp_xbar_demux_002_src0_channel;                                                                        // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                          // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                    // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                          // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                                  // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [83:0] rsp_xbar_demux_002_src1_data;                                                                           // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [25:0] rsp_xbar_demux_002_src1_channel;                                                                        // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                          // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                    // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                          // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                                  // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [83:0] rsp_xbar_demux_003_src0_data;                                                                           // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire  [25:0] rsp_xbar_demux_003_src0_channel;                                                                        // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                          // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                                    // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                          // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                                  // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [83:0] rsp_xbar_demux_003_src1_data;                                                                           // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire  [25:0] rsp_xbar_demux_003_src1_channel;                                                                        // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                          // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                    // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                          // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                                  // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [83:0] rsp_xbar_demux_004_src0_data;                                                                           // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire  [25:0] rsp_xbar_demux_004_src0_channel;                                                                        // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                          // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                    // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                          // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                                  // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [83:0] rsp_xbar_demux_005_src0_data;                                                                           // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [25:0] rsp_xbar_demux_005_src0_channel;                                                                        // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                          // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                    // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                          // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                                  // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [83:0] rsp_xbar_demux_006_src0_data;                                                                           // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [25:0] rsp_xbar_demux_006_src0_channel;                                                                        // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                          // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                    // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                          // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                                  // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [83:0] rsp_xbar_demux_007_src0_data;                                                                           // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [25:0] rsp_xbar_demux_007_src0_channel;                                                                        // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                          // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                    // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                          // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                                  // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [83:0] rsp_xbar_demux_008_src0_data;                                                                           // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire  [25:0] rsp_xbar_demux_008_src0_channel;                                                                        // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                          // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                    // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                          // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                                  // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [83:0] rsp_xbar_demux_009_src0_data;                                                                           // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire  [25:0] rsp_xbar_demux_009_src0_channel;                                                                        // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                          // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                    // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                          // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                                  // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [83:0] rsp_xbar_demux_010_src0_data;                                                                           // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire  [25:0] rsp_xbar_demux_010_src0_channel;                                                                        // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                          // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                                    // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                          // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                                  // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [83:0] rsp_xbar_demux_011_src0_data;                                                                           // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire  [25:0] rsp_xbar_demux_011_src0_channel;                                                                        // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                          // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                                    // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                          // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                                  // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [83:0] rsp_xbar_demux_012_src0_data;                                                                           // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire  [25:0] rsp_xbar_demux_012_src0_channel;                                                                        // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                          // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                                    // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                          // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                                  // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [83:0] rsp_xbar_demux_013_src0_data;                                                                           // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire  [25:0] rsp_xbar_demux_013_src0_channel;                                                                        // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                          // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_014_src0_endofpacket;                                                                    // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire         rsp_xbar_demux_014_src0_valid;                                                                          // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire         rsp_xbar_demux_014_src0_startofpacket;                                                                  // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [83:0] rsp_xbar_demux_014_src0_data;                                                                           // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire  [25:0] rsp_xbar_demux_014_src0_channel;                                                                        // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire         rsp_xbar_demux_014_src0_ready;                                                                          // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire         rsp_xbar_demux_015_src0_endofpacket;                                                                    // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire         rsp_xbar_demux_015_src0_valid;                                                                          // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire         rsp_xbar_demux_015_src0_startofpacket;                                                                  // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [83:0] rsp_xbar_demux_015_src0_data;                                                                           // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire  [25:0] rsp_xbar_demux_015_src0_channel;                                                                        // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire         rsp_xbar_demux_015_src0_ready;                                                                          // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire         rsp_xbar_demux_016_src0_endofpacket;                                                                    // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire         rsp_xbar_demux_016_src0_valid;                                                                          // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire         rsp_xbar_demux_016_src0_startofpacket;                                                                  // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [83:0] rsp_xbar_demux_016_src0_data;                                                                           // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire  [25:0] rsp_xbar_demux_016_src0_channel;                                                                        // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire         rsp_xbar_demux_016_src0_ready;                                                                          // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire         rsp_xbar_demux_017_src0_endofpacket;                                                                    // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire         rsp_xbar_demux_017_src0_valid;                                                                          // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire         rsp_xbar_demux_017_src0_startofpacket;                                                                  // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [83:0] rsp_xbar_demux_017_src0_data;                                                                           // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire  [25:0] rsp_xbar_demux_017_src0_channel;                                                                        // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire         rsp_xbar_demux_017_src0_ready;                                                                          // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire         rsp_xbar_demux_018_src0_endofpacket;                                                                    // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire         rsp_xbar_demux_018_src0_valid;                                                                          // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire         rsp_xbar_demux_018_src0_startofpacket;                                                                  // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [83:0] rsp_xbar_demux_018_src0_data;                                                                           // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire  [25:0] rsp_xbar_demux_018_src0_channel;                                                                        // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire         rsp_xbar_demux_018_src0_ready;                                                                          // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire         rsp_xbar_demux_019_src0_endofpacket;                                                                    // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire         rsp_xbar_demux_019_src0_valid;                                                                          // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	wire         rsp_xbar_demux_019_src0_startofpacket;                                                                  // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [83:0] rsp_xbar_demux_019_src0_data;                                                                           // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	wire  [25:0] rsp_xbar_demux_019_src0_channel;                                                                        // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	wire         rsp_xbar_demux_019_src0_ready;                                                                          // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire         rsp_xbar_demux_020_src0_endofpacket;                                                                    // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire         rsp_xbar_demux_020_src0_valid;                                                                          // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	wire         rsp_xbar_demux_020_src0_startofpacket;                                                                  // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [83:0] rsp_xbar_demux_020_src0_data;                                                                           // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	wire  [25:0] rsp_xbar_demux_020_src0_channel;                                                                        // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	wire         rsp_xbar_demux_020_src0_ready;                                                                          // rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire         rsp_xbar_demux_021_src0_endofpacket;                                                                    // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire         rsp_xbar_demux_021_src0_valid;                                                                          // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	wire         rsp_xbar_demux_021_src0_startofpacket;                                                                  // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [83:0] rsp_xbar_demux_021_src0_data;                                                                           // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	wire  [25:0] rsp_xbar_demux_021_src0_channel;                                                                        // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	wire         rsp_xbar_demux_021_src0_ready;                                                                          // rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire         rsp_xbar_demux_022_src0_endofpacket;                                                                    // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	wire         rsp_xbar_demux_022_src0_valid;                                                                          // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	wire         rsp_xbar_demux_022_src0_startofpacket;                                                                  // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	wire  [83:0] rsp_xbar_demux_022_src0_data;                                                                           // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	wire  [25:0] rsp_xbar_demux_022_src0_channel;                                                                        // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	wire         rsp_xbar_demux_022_src0_ready;                                                                          // rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	wire         rsp_xbar_demux_023_src0_endofpacket;                                                                    // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_001:sink23_endofpacket
	wire         rsp_xbar_demux_023_src0_valid;                                                                          // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_001:sink23_valid
	wire         rsp_xbar_demux_023_src0_startofpacket;                                                                  // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_001:sink23_startofpacket
	wire  [83:0] rsp_xbar_demux_023_src0_data;                                                                           // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_001:sink23_data
	wire  [25:0] rsp_xbar_demux_023_src0_channel;                                                                        // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_001:sink23_channel
	wire         rsp_xbar_demux_023_src0_ready;                                                                          // rsp_xbar_mux_001:sink23_ready -> rsp_xbar_demux_023:src0_ready
	wire         rsp_xbar_demux_024_src0_endofpacket;                                                                    // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_001:sink24_endofpacket
	wire         rsp_xbar_demux_024_src0_valid;                                                                          // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_001:sink24_valid
	wire         rsp_xbar_demux_024_src0_startofpacket;                                                                  // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_001:sink24_startofpacket
	wire  [83:0] rsp_xbar_demux_024_src0_data;                                                                           // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_001:sink24_data
	wire  [25:0] rsp_xbar_demux_024_src0_channel;                                                                        // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_001:sink24_channel
	wire         rsp_xbar_demux_024_src0_ready;                                                                          // rsp_xbar_mux_001:sink24_ready -> rsp_xbar_demux_024:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                            // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                          // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [83:0] limiter_cmd_src_data;                                                                                   // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [25:0] limiter_cmd_src_channel;                                                                                // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                                  // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                           // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                                 // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                         // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [83:0] rsp_xbar_mux_src_data;                                                                                  // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [25:0] rsp_xbar_mux_src_channel;                                                                               // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                                 // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                        // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                              // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                      // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [83:0] addr_router_001_src_data;                                                                               // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire  [25:0] addr_router_001_src_channel;                                                                            // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                              // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                       // rsp_xbar_mux_001:src_endofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                             // rsp_xbar_mux_001:src_valid -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                     // rsp_xbar_mux_001:src_startofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [83:0] rsp_xbar_mux_001_src_data;                                                                              // rsp_xbar_mux_001:src_data -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [25:0] rsp_xbar_mux_001_src_channel;                                                                           // rsp_xbar_mux_001:src_channel -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                             // cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                           // cmd_xbar_mux:src_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                                 // cmd_xbar_mux:src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                         // cmd_xbar_mux:src_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_mux_src_data;                                                                                  // cmd_xbar_mux:src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_mux_src_channel;                                                                               // cmd_xbar_mux:src_channel -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                              // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                    // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                            // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [83:0] id_router_src_data;                                                                                     // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [25:0] id_router_src_channel;                                                                                  // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                    // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                       // cmd_xbar_mux_002:src_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                             // cmd_xbar_mux_002:src_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                     // cmd_xbar_mux_002:src_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_mux_002_src_data;                                                                              // cmd_xbar_mux_002:src_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] cmd_xbar_mux_002_src_channel;                                                                           // cmd_xbar_mux_002:src_channel -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                             // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                          // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                                // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                        // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [83:0] id_router_002_src_data;                                                                                 // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [25:0] id_router_002_src_channel;                                                                              // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                                // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                          // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                                // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                        // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [83:0] id_router_004_src_data;                                                                                 // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [25:0] id_router_004_src_channel;                                                                              // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                                // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                          // uart_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                          // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                                // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                        // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [83:0] id_router_005_src_data;                                                                                 // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [25:0] id_router_005_src_channel;                                                                              // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                                // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                          // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                                // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                        // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [83:0] id_router_006_src_data;                                                                                 // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [25:0] id_router_006_src_channel;                                                                              // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                                // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                          // timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                          // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                                // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                        // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [83:0] id_router_007_src_data;                                                                                 // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [25:0] id_router_007_src_channel;                                                                              // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                                // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                          // lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                          // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                                // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                        // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [83:0] id_router_008_src_data;                                                                                 // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [25:0] id_router_008_src_channel;                                                                              // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                                // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_demux_001_src9_ready;                                                                          // ledr_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire         id_router_009_src_endofpacket;                                                                          // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                                // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                        // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [83:0] id_router_009_src_data;                                                                                 // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [25:0] id_router_009_src_channel;                                                                              // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                                // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_demux_001_src10_ready;                                                                         // ledg_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire         id_router_010_src_endofpacket;                                                                          // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                                // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                        // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [83:0] id_router_010_src_data;                                                                                 // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [25:0] id_router_010_src_channel;                                                                              // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                                // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_demux_001_src11_ready;                                                                         // button_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire         id_router_011_src_endofpacket;                                                                          // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                                // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                        // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [83:0] id_router_011_src_data;                                                                                 // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [25:0] id_router_011_src_channel;                                                                              // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                                // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_demux_001_src12_ready;                                                                         // switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire         id_router_012_src_endofpacket;                                                                          // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                                // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                        // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [83:0] id_router_012_src_data;                                                                                 // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [25:0] id_router_012_src_channel;                                                                              // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                                // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_demux_001_src13_ready;                                                                         // SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire         id_router_013_src_endofpacket;                                                                          // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                                // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                        // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [83:0] id_router_013_src_data;                                                                                 // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire  [25:0] id_router_013_src_channel;                                                                              // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                                // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire         cmd_xbar_demux_001_src14_ready;                                                                         // SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire         id_router_014_src_endofpacket;                                                                          // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire         id_router_014_src_valid;                                                                                // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire         id_router_014_src_startofpacket;                                                                        // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [83:0] id_router_014_src_data;                                                                                 // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire  [25:0] id_router_014_src_channel;                                                                              // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire         id_router_014_src_ready;                                                                                // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire         cmd_xbar_demux_001_src15_ready;                                                                         // SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire         id_router_015_src_endofpacket;                                                                          // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire         id_router_015_src_valid;                                                                                // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire         id_router_015_src_startofpacket;                                                                        // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [83:0] id_router_015_src_data;                                                                                 // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire  [25:0] id_router_015_src_channel;                                                                              // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire         id_router_015_src_ready;                                                                                // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire         cmd_xbar_demux_001_src16_ready;                                                                         // ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire         id_router_016_src_endofpacket;                                                                          // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire         id_router_016_src_valid;                                                                                // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire         id_router_016_src_startofpacket;                                                                        // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [83:0] id_router_016_src_data;                                                                                 // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire  [25:0] id_router_016_src_channel;                                                                              // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire         id_router_016_src_ready;                                                                                // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire         cmd_xbar_demux_001_src17_ready;                                                                         // ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire         id_router_017_src_endofpacket;                                                                          // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire         id_router_017_src_valid;                                                                                // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire         id_router_017_src_startofpacket;                                                                        // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [83:0] id_router_017_src_data;                                                                                 // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire  [25:0] id_router_017_src_channel;                                                                              // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire         id_router_017_src_ready;                                                                                // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire         cmd_xbar_demux_001_src18_ready;                                                                         // VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	wire         id_router_018_src_endofpacket;                                                                          // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire         id_router_018_src_valid;                                                                                // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire         id_router_018_src_startofpacket;                                                                        // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [83:0] id_router_018_src_data;                                                                                 // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire  [25:0] id_router_018_src_channel;                                                                              // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire         id_router_018_src_ready;                                                                                // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire         cmd_xbar_demux_001_src19_ready;                                                                         // DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	wire         id_router_019_src_endofpacket;                                                                          // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire         id_router_019_src_valid;                                                                                // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire         id_router_019_src_startofpacket;                                                                        // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [83:0] id_router_019_src_data;                                                                                 // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire  [25:0] id_router_019_src_channel;                                                                              // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire         id_router_019_src_ready;                                                                                // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire         cmd_xbar_demux_001_src20_ready;                                                                         // seg7_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	wire         id_router_020_src_endofpacket;                                                                          // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire         id_router_020_src_valid;                                                                                // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire         id_router_020_src_startofpacket;                                                                        // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [83:0] id_router_020_src_data;                                                                                 // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire  [25:0] id_router_020_src_channel;                                                                              // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire         id_router_020_src_ready;                                                                                // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire         cmd_xbar_demux_001_src22_ready;                                                                         // i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src22_ready
	wire         id_router_022_src_endofpacket;                                                                          // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire         id_router_022_src_valid;                                                                                // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire         id_router_022_src_startofpacket;                                                                        // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [83:0] id_router_022_src_data;                                                                                 // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire  [25:0] id_router_022_src_channel;                                                                              // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire         id_router_022_src_ready;                                                                                // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire         cmd_xbar_demux_001_src23_ready;                                                                         // i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src23_ready
	wire         id_router_023_src_endofpacket;                                                                          // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire         id_router_023_src_valid;                                                                                // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire         id_router_023_src_startofpacket;                                                                        // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [83:0] id_router_023_src_data;                                                                                 // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire  [25:0] id_router_023_src_channel;                                                                              // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire         id_router_023_src_ready;                                                                                // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire         cmd_xbar_demux_001_src24_ready;                                                                         // sd_wp_n_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src24_ready
	wire         id_router_024_src_endofpacket;                                                                          // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire         id_router_024_src_valid;                                                                                // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire         id_router_024_src_startofpacket;                                                                        // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [83:0] id_router_024_src_data;                                                                                 // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire  [25:0] id_router_024_src_channel;                                                                              // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire         id_router_024_src_ready;                                                                                // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire         crosser_out_ready;                                                                                      // audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire         id_router_025_src_endofpacket;                                                                          // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire         id_router_025_src_valid;                                                                                // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire         id_router_025_src_startofpacket;                                                                        // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire  [83:0] id_router_025_src_data;                                                                                 // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire  [25:0] id_router_025_src_channel;                                                                              // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire         id_router_025_src_ready;                                                                                // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                       // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                             // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                     // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [83:0] cmd_xbar_mux_001_src_data;                                                                              // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire  [25:0] cmd_xbar_mux_001_src_channel;                                                                           // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                             // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire         width_adapter_src_endofpacket;                                                                          // width_adapter:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                                // width_adapter:out_valid -> burst_adapter_001:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                        // width_adapter:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [65:0] width_adapter_src_data;                                                                                 // width_adapter:out_data -> burst_adapter_001:sink0_data
	wire         width_adapter_src_ready;                                                                                // burst_adapter_001:sink0_ready -> width_adapter:out_ready
	wire  [25:0] width_adapter_src_channel;                                                                              // width_adapter:out_channel -> burst_adapter_001:sink0_channel
	wire         id_router_001_src_endofpacket;                                                                          // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_001_src_valid;                                                                                // id_router_001:src_valid -> width_adapter_001:in_valid
	wire         id_router_001_src_startofpacket;                                                                        // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [65:0] id_router_001_src_data;                                                                                 // id_router_001:src_data -> width_adapter_001:in_data
	wire  [25:0] id_router_001_src_channel;                                                                              // id_router_001:src_channel -> width_adapter_001:in_channel
	wire         id_router_001_src_ready;                                                                                // width_adapter_001:in_ready -> id_router_001:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                      // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                            // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                                    // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [83:0] width_adapter_001_src_data;                                                                             // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire         width_adapter_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire  [25:0] width_adapter_001_src_channel;                                                                          // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                       // cmd_xbar_mux_003:src_endofpacket -> width_adapter_002:in_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                             // cmd_xbar_mux_003:src_valid -> width_adapter_002:in_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                                     // cmd_xbar_mux_003:src_startofpacket -> width_adapter_002:in_startofpacket
	wire  [83:0] cmd_xbar_mux_003_src_data;                                                                              // cmd_xbar_mux_003:src_data -> width_adapter_002:in_data
	wire  [25:0] cmd_xbar_mux_003_src_channel;                                                                           // cmd_xbar_mux_003:src_channel -> width_adapter_002:in_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                             // width_adapter_002:in_ready -> cmd_xbar_mux_003:src_ready
	wire         width_adapter_002_src_endofpacket;                                                                      // width_adapter_002:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_002_src_valid;                                                                            // width_adapter_002:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_002_src_startofpacket;                                                                    // width_adapter_002:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [56:0] width_adapter_002_src_data;                                                                             // width_adapter_002:out_data -> burst_adapter:sink0_data
	wire         width_adapter_002_src_ready;                                                                            // burst_adapter:sink0_ready -> width_adapter_002:out_ready
	wire  [25:0] width_adapter_002_src_channel;                                                                          // width_adapter_002:out_channel -> burst_adapter:sink0_channel
	wire         id_router_003_src_endofpacket;                                                                          // id_router_003:src_endofpacket -> width_adapter_003:in_endofpacket
	wire         id_router_003_src_valid;                                                                                // id_router_003:src_valid -> width_adapter_003:in_valid
	wire         id_router_003_src_startofpacket;                                                                        // id_router_003:src_startofpacket -> width_adapter_003:in_startofpacket
	wire  [56:0] id_router_003_src_data;                                                                                 // id_router_003:src_data -> width_adapter_003:in_data
	wire  [25:0] id_router_003_src_channel;                                                                              // id_router_003:src_channel -> width_adapter_003:in_channel
	wire         id_router_003_src_ready;                                                                                // width_adapter_003:in_ready -> id_router_003:src_ready
	wire         width_adapter_003_src_endofpacket;                                                                      // width_adapter_003:out_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         width_adapter_003_src_valid;                                                                            // width_adapter_003:out_valid -> rsp_xbar_demux_003:sink_valid
	wire         width_adapter_003_src_startofpacket;                                                                    // width_adapter_003:out_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [83:0] width_adapter_003_src_data;                                                                             // width_adapter_003:out_data -> rsp_xbar_demux_003:sink_data
	wire         width_adapter_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> width_adapter_003:out_ready
	wire  [25:0] width_adapter_003_src_channel;                                                                          // width_adapter_003:out_channel -> rsp_xbar_demux_003:sink_channel
	wire         cmd_xbar_demux_001_src21_ready;                                                                         // width_adapter_004:in_ready -> cmd_xbar_demux_001:src21_ready
	wire         width_adapter_004_src_endofpacket;                                                                      // width_adapter_004:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire         width_adapter_004_src_valid;                                                                            // width_adapter_004:out_valid -> burst_adapter_002:sink0_valid
	wire         width_adapter_004_src_startofpacket;                                                                    // width_adapter_004:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire  [65:0] width_adapter_004_src_data;                                                                             // width_adapter_004:out_data -> burst_adapter_002:sink0_data
	wire         width_adapter_004_src_ready;                                                                            // burst_adapter_002:sink0_ready -> width_adapter_004:out_ready
	wire  [25:0] width_adapter_004_src_channel;                                                                          // width_adapter_004:out_channel -> burst_adapter_002:sink0_channel
	wire         id_router_021_src_endofpacket;                                                                          // id_router_021:src_endofpacket -> width_adapter_005:in_endofpacket
	wire         id_router_021_src_valid;                                                                                // id_router_021:src_valid -> width_adapter_005:in_valid
	wire         id_router_021_src_startofpacket;                                                                        // id_router_021:src_startofpacket -> width_adapter_005:in_startofpacket
	wire  [65:0] id_router_021_src_data;                                                                                 // id_router_021:src_data -> width_adapter_005:in_data
	wire  [25:0] id_router_021_src_channel;                                                                              // id_router_021:src_channel -> width_adapter_005:in_channel
	wire         id_router_021_src_ready;                                                                                // width_adapter_005:in_ready -> id_router_021:src_ready
	wire         width_adapter_005_src_endofpacket;                                                                      // width_adapter_005:out_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire         width_adapter_005_src_valid;                                                                            // width_adapter_005:out_valid -> rsp_xbar_demux_021:sink_valid
	wire         width_adapter_005_src_startofpacket;                                                                    // width_adapter_005:out_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [83:0] width_adapter_005_src_data;                                                                             // width_adapter_005:out_data -> rsp_xbar_demux_021:sink_data
	wire         width_adapter_005_src_ready;                                                                            // rsp_xbar_demux_021:sink_ready -> width_adapter_005:out_ready
	wire  [25:0] width_adapter_005_src_channel;                                                                          // width_adapter_005:out_channel -> rsp_xbar_demux_021:sink_channel
	wire         crosser_out_endofpacket;                                                                                // crosser:out_endofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_out_valid;                                                                                      // crosser:out_valid -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_out_startofpacket;                                                                              // crosser:out_startofpacket -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] crosser_out_data;                                                                                       // crosser:out_data -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [25:0] crosser_out_channel;                                                                                    // crosser:out_channel -> audio_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src25_endofpacket;                                                                   // cmd_xbar_demux_001:src25_endofpacket -> crosser:in_endofpacket
	wire         cmd_xbar_demux_001_src25_valid;                                                                         // cmd_xbar_demux_001:src25_valid -> crosser:in_valid
	wire         cmd_xbar_demux_001_src25_startofpacket;                                                                 // cmd_xbar_demux_001:src25_startofpacket -> crosser:in_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src25_data;                                                                          // cmd_xbar_demux_001:src25_data -> crosser:in_data
	wire  [25:0] cmd_xbar_demux_001_src25_channel;                                                                       // cmd_xbar_demux_001:src25_channel -> crosser:in_channel
	wire         cmd_xbar_demux_001_src25_ready;                                                                         // crosser:in_ready -> cmd_xbar_demux_001:src25_ready
	wire         crosser_001_out_endofpacket;                                                                            // crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink25_endofpacket
	wire         crosser_001_out_valid;                                                                                  // crosser_001:out_valid -> rsp_xbar_mux_001:sink25_valid
	wire         crosser_001_out_startofpacket;                                                                          // crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink25_startofpacket
	wire  [83:0] crosser_001_out_data;                                                                                   // crosser_001:out_data -> rsp_xbar_mux_001:sink25_data
	wire  [25:0] crosser_001_out_channel;                                                                                // crosser_001:out_channel -> rsp_xbar_mux_001:sink25_channel
	wire         crosser_001_out_ready;                                                                                  // rsp_xbar_mux_001:sink25_ready -> crosser_001:out_ready
	wire         rsp_xbar_demux_025_src0_endofpacket;                                                                    // rsp_xbar_demux_025:src0_endofpacket -> crosser_001:in_endofpacket
	wire         rsp_xbar_demux_025_src0_valid;                                                                          // rsp_xbar_demux_025:src0_valid -> crosser_001:in_valid
	wire         rsp_xbar_demux_025_src0_startofpacket;                                                                  // rsp_xbar_demux_025:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [83:0] rsp_xbar_demux_025_src0_data;                                                                           // rsp_xbar_demux_025:src0_data -> crosser_001:in_data
	wire  [25:0] rsp_xbar_demux_025_src0_channel;                                                                        // rsp_xbar_demux_025:src0_channel -> crosser_001:in_channel
	wire         rsp_xbar_demux_025_src0_ready;                                                                          // crosser_001:in_ready -> rsp_xbar_demux_025:src0_ready
	wire  [25:0] limiter_cmd_valid_data;                                                                                 // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                               // epcs_controller:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                               // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                               // uart_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                               // timer_0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                                               // timer_1:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                                               // button_pio:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                                                               // DM9000A:oINT -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                                                               // ISP1362:avs_dc_irq_n_oINT0_N -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                                                                               // ISP1362:avs_hc_irq_n_oINT0_N -> irq_mapper:receiver8_irq
	wire  [31:0] cpu_0_d_irq_irq;                                                                                        // irq_mapper:sender_irq -> cpu_0:d_irq

	system_0_sdram_0 sdram_0 (
		.clk            (clk),                                                     //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                         // reset.reset_n
		.az_addr        (sdram_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram_0),                                //  wire.export
		.zs_ba          (zs_ba_from_the_sdram_0),                                  //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram_0),                               //      .export
		.zs_cke         (zs_cke_from_the_sdram_0),                                 //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram_0),                                //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram_0),                           //      .export
		.zs_dqm         (zs_dqm_from_the_sdram_0),                                 //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram_0),                               //      .export
		.zs_we_n        (zs_we_n_from_the_sdram_0)                                 //      .export
	);

	system_0_epcs_controller epcs_controller (
		.clk           (clk),                                                                         //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                             //             reset.reset_n
		.address       (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address),    // epcs_control_port.address
		.chipselect    (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect), //                  .chipselect
		.dataavailable (),                                                                            //                  .dataavailable
		.endofpacket   (),                                                                            //                  .endofpacket
		.read_n        (~epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read),      //                  .read_n
		.readdata      (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata),   //                  .readdata
		.readyfordata  (),                                                                            //                  .readyfordata
		.write_n       (~epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write),     //                  .write_n
		.writedata     (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver0_irq)                                                     //               irq.irq
	);

	system_0_jtag_uart_0 jtag_uart_0 (
		.clk            (clk),                                                                      //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.dataavailable  (),                                                                         //                  .dataavailable
		.readyfordata   (),                                                                         //                  .readyfordata
		.av_irq         (irq_mapper_receiver1_irq)                                                  //               irq.irq
	);

	system_0_uart_0 uart_0 (
		.clk           (clk),                                                    //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address       (uart_0_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_0_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_0_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_0_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_0_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_0_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_0_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                       //                    .dataavailable
		.readyfordata  (),                                                       //                    .readyfordata
		.rxd           (rxd_to_the_uart_0),                                      // external_connection.export
		.txd           (txd_from_the_uart_0),                                    //                    .export
		.irq           (irq_mapper_receiver2_irq)                                //                 irq.irq
	);

	system_0_timer_0 timer_0 (
		.clk        (clk),                                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                              //   irq.irq
	);

	system_0_timer_0 timer_1 (
		.clk        (clk),                                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                              //   irq.irq
	);

	system_0_lcd lcd (
		.clk           (clk),                                                            //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                //         reset.reset_n
		.address       (lcd_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (lcd_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.read          (lcd_control_slave_translator_avalon_anti_slave_0_read),          //              .read
		.readdata      (lcd_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (lcd_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (lcd_control_slave_translator_avalon_anti_slave_0_writedata),     //              .writedata
		.LCD_data      (LCD_data_to_and_from_the_lcd_16207_0),                           //      external.export
		.LCD_E         (LCD_E_from_the_lcd_16207_0),                                     //              .export
		.LCD_RS        (LCD_RS_from_the_lcd_16207_0),                                    //              .export
		.LCD_RW        (LCD_RW_from_the_lcd_16207_0)                                     //              .export
	);

	system_0_ledr ledr (
		.clk        (clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledr_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledr_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledr_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledr_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledr_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led_red)                          // external_connection.export
	);

	system_0_ledg ledg (
		.clk        (clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledg_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledg_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledg_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledg_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledg_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led_green)                        // external_connection.export
	);

	system_0_button_pio button_pio (
		.clk        (clk),                                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (button_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~button_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (button_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (button_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (button_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (in_port_to_the_button_pio),                               // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                                 //                 irq.irq
	);

	system_0_switch_pio switch_pio (
		.clk      (clk),                                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (switch_pio_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switch_pio_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (in_port_to_the_switch_pio)                              // external_connection.export
	);

	system_0_SD_DAT sd_dat (
		.clk        (clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (sd_dat_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sd_dat_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sd_dat_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sd_dat_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sd_dat_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (bidir_port_to_and_from_the_SD_DAT)                    // external_connection.export
	);

	system_0_SD_CMD sd_cmd (
		.clk        (clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (sd_cmd_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sd_cmd_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sd_cmd_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sd_cmd_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sd_cmd_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (bidir_port_to_and_from_the_SD_CMD)                    // external_connection.export
	);

	system_0_SD_CLK sd_clk (
		.clk        (clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (sd_clk_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sd_clk_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sd_clk_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sd_clk_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sd_clk_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_SD_CLK)                             // external_connection.export
	);

	ISP1362_IF isp1362 (
		.avs_hc_clk_iCLK           (clk),                                                   //    hc_clock.clk
		.avs_hc_reset_n_iRST_N     (~rst_controller_001_reset_out_reset),                   //  hc_reset_n.reset_n
		.avs_hc_writedata_iDATA    (isp1362_hc_translator_avalon_anti_slave_0_writedata),   //          hc.writedata
		.avs_hc_readdata_oDATA     (isp1362_hc_translator_avalon_anti_slave_0_readdata),    //            .readdata
		.avs_hc_address_iADDR      (isp1362_hc_translator_avalon_anti_slave_0_address),     //            .address
		.avs_hc_read_n_iRD_N       (~isp1362_hc_translator_avalon_anti_slave_0_read),       //            .read_n
		.avs_hc_write_n_iWR_N      (~isp1362_hc_translator_avalon_anti_slave_0_write),      //            .write_n
		.avs_hc_chipselect_n_iCS_N (~isp1362_hc_translator_avalon_anti_slave_0_chipselect), //            .chipselect_n
		.avs_hc_irq_n_oINT0_N      (irq_mapper_receiver8_irq),                              //      hc_irq.irq_n
		.avs_dc_clk_iCLK           (clk),                                                   //    dc_clock.clk
		.avs_dc_reset_n_iRST_N     (~rst_controller_001_reset_out_reset),                   //  dc_reset_n.reset_n
		.avs_dc_writedata_iDATA    (isp1362_dc_translator_avalon_anti_slave_0_writedata),   //          dc.writedata
		.avs_dc_readdata_oDATA     (isp1362_dc_translator_avalon_anti_slave_0_readdata),    //            .readdata
		.avs_dc_address_iADDR      (isp1362_dc_translator_avalon_anti_slave_0_address),     //            .address
		.avs_dc_read_n_iRD_N       (~isp1362_dc_translator_avalon_anti_slave_0_read),       //            .read_n
		.avs_dc_write_n_iWR_N      (~isp1362_dc_translator_avalon_anti_slave_0_write),      //            .write_n
		.avs_dc_chipselect_n_iCS_N (~isp1362_dc_translator_avalon_anti_slave_0_chipselect), //            .chipselect_n
		.avs_dc_irq_n_oINT0_N      (irq_mapper_receiver7_irq),                              //      dc_irq.irq_n
		.USB_DATA                  (ISP1362_conduit_end_DATA),                              // conduit_end.export
		.USB_ADDR                  (ISP1362_conduit_end_ADDR),                              //            .export
		.USB_RD_N                  (ISP1362_conduit_end_RD_N),                              //            .export
		.USB_WR_N                  (ISP1362_conduit_end_WR_N),                              //            .export
		.USB_CS_N                  (ISP1362_conduit_end_CS_N),                              //            .export
		.USB_RST_N                 (ISP1362_conduit_end_RST_N),                             //            .export
		.USB_INT0                  (ISP1362_conduit_end_INT0),                              //            .export
		.USB_INT1                  (ISP1362_conduit_end_INT1)                               //            .export
	);

	system_0_cpu_0 cpu_0 (
		.clk                                   (clk),                                                                  //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (cpu_0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_0_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_0_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_0_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_0_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	system_0_tri_state_bridge_0_bridge_0 tri_state_bridge_0_bridge_0 (
		.clk                               (clk),                                                                //   clk.clk
		.reset                             (rst_controller_reset_out_reset),                                     // reset.reset
		.request                           (tri_state_bridge_0_pinsharer_0_tcm_request),                         //   tcs.request
		.grant                             (tri_state_bridge_0_pinsharer_0_tcm_grant),                           //      .grant
		.tcs_tri_state_bridge_0_data       (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out),     //      .tri_state_bridge_0_data_out
		.tcs_tri_state_bridge_0_data_outen (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen),   //      .tri_state_bridge_0_data_outen
		.tcs_tri_state_bridge_0_data_in    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in),      //      .tri_state_bridge_0_data_in
		.tcs_tri_state_bridge_0_readn      (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out),    //      .tri_state_bridge_0_readn_out
		.tcs_write_n_to_the_cfi_flash_0    (tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out),  //      .write_n_to_the_cfi_flash_0_out
		.tcs_tri_state_bridge_0_address    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out),  //      .tri_state_bridge_0_address_out
		.tcs_select_n_to_the_cfi_flash_0   (tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out), //      .select_n_to_the_cfi_flash_0_out
		.tri_state_bridge_0_data           (tri_state_bridge_0_data),                                            //   out.tri_state_bridge_0_data
		.tri_state_bridge_0_readn          (tri_state_bridge_0_readn),                                           //      .tri_state_bridge_0_readn
		.write_n_to_the_cfi_flash_0        (write_n_to_the_cfi_flash_0),                                         //      .write_n_to_the_cfi_flash_0
		.tri_state_bridge_0_address        (tri_state_bridge_0_address),                                         //      .tri_state_bridge_0_address
		.select_n_to_the_cfi_flash_0       (select_n_to_the_cfi_flash_0)                                         //      .select_n_to_the_cfi_flash_0
	);

	system_0_tri_state_bridge_0_pinSharer_0 tri_state_bridge_0_pinsharer_0 (
		.clk_clk                       (clk),                                                                //   clk.clk
		.reset_reset                   (rst_controller_reset_out_reset),                                     // reset.reset
		.request                       (tri_state_bridge_0_pinsharer_0_tcm_request),                         //   tcm.request
		.grant                         (tri_state_bridge_0_pinsharer_0_tcm_grant),                           //      .grant
		.tri_state_bridge_0_address    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out),  //      .tri_state_bridge_0_address_out
		.tri_state_bridge_0_readn      (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out),    //      .tri_state_bridge_0_readn_out
		.write_n_to_the_cfi_flash_0    (tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out),  //      .write_n_to_the_cfi_flash_0_out
		.tri_state_bridge_0_data       (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out),     //      .tri_state_bridge_0_data_out
		.tri_state_bridge_0_data_in    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in),      //      .tri_state_bridge_0_data_in
		.tri_state_bridge_0_data_outen (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen),   //      .tri_state_bridge_0_data_outen
		.select_n_to_the_cfi_flash_0   (tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out), //      .select_n_to_the_cfi_flash_0_out
		.tcs0_request                  (cfi_flash_0_tcm_request),                                            //  tcs0.request
		.tcs0_grant                    (cfi_flash_0_tcm_grant),                                              //      .grant
		.tcs0_address_out              (cfi_flash_0_tcm_address_out),                                        //      .address_out
		.tcs0_read_n_out               (cfi_flash_0_tcm_read_n_out),                                         //      .read_n_out
		.tcs0_write_n_out              (cfi_flash_0_tcm_write_n_out),                                        //      .write_n_out
		.tcs0_data_out                 (cfi_flash_0_tcm_data_out),                                           //      .data_out
		.tcs0_data_in                  (cfi_flash_0_tcm_data_in),                                            //      .data_in
		.tcs0_data_outen               (cfi_flash_0_tcm_data_outen),                                         //      .data_outen
		.tcs0_chipselect_n_out         (cfi_flash_0_tcm_chipselect_n_out)                                    //      .chipselect_n_out
	);

	system_0_cfi_flash_0 #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (40),
		.TCM_DATA_HOLD                  (40),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) cfi_flash_0 (
		.clk_clk              (clk),                                                          //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                               // reset.reset
		.uas_address          (cfi_flash_0_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (cfi_flash_0_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (cfi_flash_0_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (cfi_flash_0_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (cfi_flash_0_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (cfi_flash_0_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (cfi_flash_0_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (cfi_flash_0_tcm_request),                                      //      .request
		.tcm_grant            (cfi_flash_0_tcm_grant),                                        //      .grant
		.tcm_address_out      (cfi_flash_0_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (cfi_flash_0_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (cfi_flash_0_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (cfi_flash_0_tcm_data_in)                                       //      .data_in
	);

	VGA_NIOS_CTRL #(
		.RAM_SIZE (307200)
	) vga_0 (
		.iCLK      (clk),                                                            //                   clk.clk
		.VGA_R     (vga_0_avalon_slave_0_export_VGA_R),                              // avalon_slave_0_export.export
		.VGA_G     (vga_0_avalon_slave_0_export_VGA_G),                              //                      .export
		.VGA_B     (vga_0_avalon_slave_0_export_VGA_B),                              //                      .export
		.VGA_HS    (vga_0_avalon_slave_0_export_VGA_HS),                             //                      .export
		.VGA_VS    (vga_0_avalon_slave_0_export_VGA_VS),                             //                      .export
		.VGA_SYNC  (vga_0_avalon_slave_0_export_VGA_SYNC),                           //                      .export
		.VGA_BLANK (vga_0_avalon_slave_0_export_VGA_BLANK),                          //                      .export
		.VGA_CLK   (vga_0_avalon_slave_0_export_VGA_CLK),                            //                      .export
		.iCLK_25   (vga_0_avalon_slave_0_export_iCLK_25),                            //                      .export
		.oDATA     (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //        avalon_slave_0.readdata
		.iDATA     (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //                      .writedata
		.iADDR     (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //                      .address
		.iWR       (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //                      .write
		.iRD       (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //                      .read
		.iCS       (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //                      .chipselect
		.iRST_N    (~rst_controller_001_reset_out_reset)                             //               reset_n.reset_n
	);

	DM9000A_IF dm9000a (
		.iCLK       (clk),                                                               //                   clk.clk
		.iOSC_50    (dm9000a_avalon_slave_0_export_iOSC_50),                             // avalon_slave_0_export.export
		.ENET_DATA  (dm9000a_avalon_slave_0_export_ENET_DATA),                           //                      .export
		.ENET_CMD   (dm9000a_avalon_slave_0_export_ENET_CMD),                            //                      .export
		.ENET_RD_N  (dm9000a_avalon_slave_0_export_ENET_RD_N),                           //                      .export
		.ENET_WR_N  (dm9000a_avalon_slave_0_export_ENET_WR_N),                           //                      .export
		.ENET_CS_N  (dm9000a_avalon_slave_0_export_ENET_CS_N),                           //                      .export
		.ENET_RST_N (dm9000a_avalon_slave_0_export_ENET_RST_N),                          //                      .export
		.ENET_CLK   (dm9000a_avalon_slave_0_export_ENET_CLK),                            //                      .export
		.ENET_INT   (dm9000a_avalon_slave_0_export_ENET_INT),                            //                      .export
		.iDATA      (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //        avalon_slave_0.writedata
		.iCMD       (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address),     //                      .address
		.iRD_N      (~dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read),       //                      .read_n
		.iWR_N      (~dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write),      //                      .write_n
		.iCS_N      (~dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //                      .chipselect_n
		.oDATA      (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                      .readdata
		.oINT       (irq_mapper_receiver6_irq),                                          //    avalon_slave_0_irq.irq
		.iRST_N     (~rst_controller_001_reset_out_reset)                                //               reset_n.reset_n
	);

	SEG7_LUT_8 seg7 (
		.iCLK   (clk),                                                        //          clk.clk
		.iWR    (seg7_avalon_slave_translator_avalon_anti_slave_0_write),     // avalon_slave.write
		.iDIG   (seg7_avalon_slave_translator_avalon_anti_slave_0_writedata), //             .writedata
		.oSEG0  (seg7_display_conduit_end_oSEG0),                             //  conduit_end.export
		.oSEG1  (seg7_display_conduit_end_oSEG1),                             //             .export
		.oSEG2  (seg7_display_conduit_end_oSEG2),                             //             .export
		.oSEG3  (seg7_display_conduit_end_oSEG3),                             //             .export
		.oSEG4  (seg7_display_conduit_end_oSEG4),                             //             .export
		.oSEG5  (seg7_display_conduit_end_oSEG5),                             //             .export
		.oSEG6  (seg7_display_conduit_end_oSEG6),                             //             .export
		.oSEG7  (seg7_display_conduit_end_oSEG7),                             //             .export
		.iRST_N (~rst_controller_001_reset_out_reset)                         //      reset_n.reset_n
	);

	SRAM_16Bit_512K sram_0 (
		.iCLK      (clk),                                                              //                   clk.clk
		.SRAM_DQ   (sram_0_avalon_slave_0_export_DQ),                                  // avalon_slave_0_export.export
		.SRAM_ADDR (sram_0_avalon_slave_0_export_ADDR),                                //                      .export
		.SRAM_UB_N (sram_0_avalon_slave_0_export_UB_N),                                //                      .export
		.SRAM_LB_N (sram_0_avalon_slave_0_export_LB_N),                                //                      .export
		.SRAM_WE_N (sram_0_avalon_slave_0_export_WE_N),                                //                      .export
		.SRAM_CE_N (sram_0_avalon_slave_0_export_CE_N),                                //                      .export
		.SRAM_OE_N (sram_0_avalon_slave_0_export_OE_N),                                //                      .export
		.iDATA     (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //        avalon_slave_0.writedata
		.oDATA     (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                      .readdata
		.iADDR     (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_address),     //                      .address
		.iWE_N     (~sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //                      .write_n
		.iOE_N     (~sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //                      .read_n
		.iCE_N     (~sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //                      .chipselect_n
		.iBE_N     (~sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //                      .byteenable_n
		.iRST_N    (~rst_controller_001_reset_out_reset)                               //               reset_n.reset_n
	);

	system_0_SD_CLK i2c_scl (
		.clk        (clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (i2c_scl_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_scl_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_scl_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_scl_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_scl_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)                    // external_connection.export
	);

	system_0_SD_CMD i2c_sda (
		.clk        (clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (i2c_sda_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~i2c_sda_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (i2c_sda_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (i2c_sda_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (i2c_sda_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)                    // external_connection.export
	);

	system_0_sd_wp_n sd_wp_n (
		.clk      (clk),                                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                //               reset.reset_n
		.address  (sd_wp_n_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (sd_wp_n_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (sd_wp_n_external_connection_export)                  // external_connection.export
	);

	AUDIO_IF audio (
		.avs_s1_address       (audio_avalon_slave_translator_avalon_anti_slave_0_address),   //     avalon_slave.address
		.avs_s1_read          (audio_avalon_slave_translator_avalon_anti_slave_0_read),      //                 .read
		.avs_s1_readdata      (audio_avalon_slave_translator_avalon_anti_slave_0_readdata),  //                 .readdata
		.avs_s1_write         (audio_avalon_slave_translator_avalon_anti_slave_0_write),     //                 .write
		.avs_s1_writedata     (audio_avalon_slave_translator_avalon_anti_slave_0_writedata), //                 .writedata
		.avs_s1_clk           (clk_audio_clk_in_clk),                                        //       clock_sink.clk
		.avs_s1_reset         (rst_controller_002_reset_out_reset),                          // clock_sink_reset.reset
		.avs_s1_export_XCK    (audio_conduit_end_XCK),                                       //      conduit_end.export
		.avs_s1_export_ADCDAT (audio_conduit_end_ADCDAT),                                    //                 .export
		.avs_s1_export_ADCLRC (audio_conduit_end_ADCLRC),                                    //                 .export
		.avs_s1_export_DACDAT (audio_conduit_end_DACDAT),                                    //                 .export
		.avs_s1_export_DACLRC (audio_conduit_end_DACLRC),                                    //                 .export
		.avs_s1_export_BCLK   (audio_conduit_end_BCLK)                                       //                 .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_0_instruction_master_translator (
		.clk                   (clk),                                                                         //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_0_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_0_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_0_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_0_data_master_translator (
		.clk                   (clk),                                                                  //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_0_data_master_read),                                               //                          .read
		.av_readdata           (cpu_0_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_0_data_master_write),                                              //                          .write
		.av_writedata          (cpu_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_0_jtag_debug_module_translator (
		.clk                   (clk),                                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_0_s1_translator (
		.clk                   (clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) epcs_controller_epcs_control_port_translator (
		.clk                   (clk),                                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                               //                    reset.reset
		.uav_address           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_byteenable         (),                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_debugaccess        (),                                                                                             //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cfi_flash_0_uas_translator (
		.clk                   (clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                             //                    reset.reset
		.uav_address           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cfi_flash_0_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cfi_flash_0_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (cfi_flash_0_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (cfi_flash_0_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_chipselect         (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (clk),                                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_0_s1_translator (
		.clk                   (clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (uart_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (uart_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (uart_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (uart_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (uart_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (uart_0_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect         (uart_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_1_s1_translator (
		.clk                   (clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (25),
		.AV_WRITE_WAIT_CYCLES           (25),
		.AV_SETUP_WAIT_CYCLES           (25),
		.AV_DATA_HOLD_CYCLES            (25)
	) lcd_control_slave_translator (
		.clk                   (clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (lcd_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (lcd_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (lcd_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (lcd_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (lcd_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (lcd_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledr_s1_translator (
		.clk                   (clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ledr_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ledr_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ledr_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ledr_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (ledr_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledg_s1_translator (
		.clk                   (clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ledg_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ledg_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ledg_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ledg_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (ledg_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_pio_s1_translator (
		.clk                   (clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (button_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (button_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (button_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (button_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (button_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch_pio_s1_translator (
		.clk                   (clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switch_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (switch_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                         //              (terminated)
		.av_read               (),                                                                         //              (terminated)
		.av_writedata          (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_dat_s1_translator (
		.clk                   (clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_dat_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_dat_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sd_dat_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_dat_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_dat_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_cmd_s1_translator (
		.clk                   (clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_cmd_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_cmd_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sd_cmd_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_cmd_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_cmd_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_clk_s1_translator (
		.clk                   (clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_clk_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_clk_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sd_clk_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_clk_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_clk_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (15),
		.AV_WRITE_WAIT_CYCLES           (15),
		.AV_SETUP_WAIT_CYCLES           (15),
		.AV_DATA_HOLD_CYCLES            (15)
	) isp1362_dc_translator (
		.clk                   (clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (isp1362_dc_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (isp1362_dc_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (isp1362_dc_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (isp1362_dc_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (isp1362_dc_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (isp1362_dc_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (5),
		.AV_WRITE_WAIT_CYCLES           (5),
		.AV_SETUP_WAIT_CYCLES           (14),
		.AV_DATA_HOLD_CYCLES            (14)
	) isp1362_hc_translator (
		.clk                   (clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (isp1362_hc_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (isp1362_hc_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (isp1362_hc_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (isp1362_hc_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (isp1362_hc_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (isp1362_hc_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (19),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (1),
		.AV_DATA_HOLD_CYCLES            (1)
	) vga_0_avalon_slave_0_translator (
		.clk                   (clk),                                                                             //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address           (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (vga_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (4),
		.AV_WRITE_WAIT_CYCLES           (4),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dm9000a_avalon_slave_0_translator (
		.clk                   (clk),                                                                               //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seg7_avalon_slave_translator (
		.clk                   (clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (seg7_avalon_slave_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (seg7_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_address            (),                                                                             //              (terminated)
		.av_read               (),                                                                             //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                         //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (2),
		.AV_WRITE_WAIT_CYCLES           (2),
		.AV_SETUP_WAIT_CYCLES           (2),
		.AV_DATA_HOLD_CYCLES            (2)
	) sram_0_avalon_slave_0_translator (
		.clk                   (clk),                                                                              //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                               //                    reset.reset
		.uav_address           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_sda_s1_translator (
		.clk                   (clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (i2c_sda_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (i2c_sda_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (i2c_sda_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (i2c_sda_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (i2c_sda_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) i2c_scl_s1_translator (
		.clk                   (clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (i2c_scl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (i2c_scl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (i2c_scl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (i2c_scl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (i2c_scl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_wp_n_s1_translator (
		.clk                   (clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_wp_n_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sd_wp_n_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                      //              (terminated)
		.av_read               (),                                                                      //              (terminated)
		.av_writedata          (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_chipselect         (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_avalon_slave_translator (
		.clk                   (clk_audio_clk_in_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                            //                    reset.reset
		.uav_address           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (audio_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (audio_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (audio_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (audio_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) lcd_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                        //                .channel
		.rf_sink_ready           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) isp1362_hc_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (isp1362_hc_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                                //                .channel
		.rf_sink_ready           (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_wp_n_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src24_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src24_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src24_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src24_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src24_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src24_channel),                                                //                .channel
		.rf_sink_ready           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switch_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                   //                .channel
		.rf_sink_ready           (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ledg_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                             //                .channel
		.rf_sink_ready           (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) i2c_sda_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src22_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src22_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src22_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src22_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src22_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src22_channel),                                                //                .channel
		.rf_sink_ready           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) button_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                   //                .channel
		.rf_sink_ready           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ledr_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                              //                .channel
		.rf_sink_ready           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) seg7_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src20_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src20_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src20_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src20_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src20_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src20_channel),                                                       //                .channel
		.rf_sink_ready           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (45),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_POSTED          (35),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.PKT_TRANS_LOCK            (38),
		.PKT_SRC_ID_H              (50),
		.PKT_SRC_ID_L              (46),
		.PKT_DEST_ID_H             (55),
		.PKT_DEST_ID_L             (51),
		.PKT_BURSTWRAP_H           (44),
		.PKT_BURSTWRAP_L           (42),
		.PKT_BYTE_CNT_H            (41),
		.PKT_BYTE_CNT_L            (39),
		.PKT_PROTECTION_H          (56),
		.PKT_PROTECTION_L          (56),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (57),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cfi_flash_0_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                          //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                          //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                           //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                    //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                        //                .channel
		.rf_sink_ready           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (58),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                 //                .channel
		.rf_sink_ready           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_cmd_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                               //                .channel
		.rf_sink_ready           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) uart_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                //                .channel
		.rf_sink_ready           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src19_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src19_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src19_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src19_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src19_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src19_channel),                                                            //                .channel
		.rf_sink_ready           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) isp1362_dc_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (isp1362_dc_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                //                .channel
		.rf_sink_ready           (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src18_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src18_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src18_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src18_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src18_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src18_channel),                                                          //                .channel
		.rf_sink_ready           (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_audio_clk_in_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                       //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                       //                .valid
		.cp_data                 (crosser_out_data),                                                                        //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                     //                .channel
		.rf_sink_ready           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_audio_clk_in_clk),                                                                    //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_audio_clk_in_clk),                                                              //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                // clk_reset.reset
		.in_data           (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_clk_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                               //                .channel
		.rf_sink_ready           (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                           //                .channel
		.rf_sink_ready           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (26),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) cpu_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk),                                                                           //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                     //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                 //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_dat_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                               //                .channel
		.rf_sink_ready           (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (26),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3)
	) cpu_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk),                                                                                  //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                 //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                              //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                        //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                          //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                 //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (54),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (59),
		.PKT_SRC_ID_L              (55),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (60),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                 //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                 //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                  //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                           //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                               //                .channel
		.rf_sink_ready           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) i2c_scl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src23_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src23_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src23_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src23_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src23_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src23_channel),                                                //                .channel
		.rf_sink_ready           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (54),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (59),
		.PKT_SRC_ID_L              (55),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (60),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (26),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                            //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                            //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                             //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                          //                .channel
		.rf_sink_ready           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	system_0_addr_router addr_router (
		.sink_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	system_0_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	system_0_id_router id_router (
		.sink_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	system_0_id_router_001 id_router_001 (
		.sink_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                               //       src.ready
		.src_valid          (id_router_001_src_valid),                                               //          .valid
		.src_data           (id_router_001_src_data),                                                //          .data
		.src_channel        (id_router_001_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router id_router_002 (
		.sink_ready         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                      //          .valid
		.src_data           (id_router_002_src_data),                                                                       //          .data
		.src_channel        (id_router_002_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                                 //          .endofpacket
	);

	system_0_id_router_003 id_router_003 (
		.sink_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                    //       src.ready
		.src_valid          (id_router_003_src_valid),                                                    //          .valid
		.src_data           (id_router_003_src_data),                                                     //          .data
		.src_channel        (id_router_003_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                               //          .endofpacket
	);

	system_0_id_router_004 id_router_004 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                  //          .valid
		.src_data           (id_router_004_src_data),                                                                   //          .data
		.src_channel        (id_router_004_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                             //          .endofpacket
	);

	system_0_id_router_004 id_router_005 (
		.sink_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                              //       src.ready
		.src_valid          (id_router_005_src_valid),                                              //          .valid
		.src_data           (id_router_005_src_data),                                               //          .data
		.src_channel        (id_router_005_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                         //          .endofpacket
	);

	system_0_id_router_004 id_router_006 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                               //       src.ready
		.src_valid          (id_router_006_src_valid),                                               //          .valid
		.src_data           (id_router_006_src_data),                                                //          .data
		.src_channel        (id_router_006_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_004 id_router_007 (
		.sink_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                               //       src.ready
		.src_valid          (id_router_007_src_valid),                                               //          .valid
		.src_data           (id_router_007_src_data),                                                //          .data
		.src_channel        (id_router_007_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_004 id_router_008 (
		.sink_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                      //       src.ready
		.src_valid          (id_router_008_src_valid),                                                      //          .valid
		.src_data           (id_router_008_src_data),                                                       //          .data
		.src_channel        (id_router_008_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                 //          .endofpacket
	);

	system_0_id_router_004 id_router_009 (
		.sink_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                            //       src.ready
		.src_valid          (id_router_009_src_valid),                                            //          .valid
		.src_data           (id_router_009_src_data),                                             //          .data
		.src_channel        (id_router_009_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                       //          .endofpacket
	);

	system_0_id_router_004 id_router_010 (
		.sink_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                            //       src.ready
		.src_valid          (id_router_010_src_valid),                                            //          .valid
		.src_data           (id_router_010_src_data),                                             //          .data
		.src_channel        (id_router_010_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                       //          .endofpacket
	);

	system_0_id_router_004 id_router_011 (
		.sink_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                  //       src.ready
		.src_valid          (id_router_011_src_valid),                                                  //          .valid
		.src_data           (id_router_011_src_data),                                                   //          .data
		.src_channel        (id_router_011_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                             //          .endofpacket
	);

	system_0_id_router_004 id_router_012 (
		.sink_ready         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                  //       src.ready
		.src_valid          (id_router_012_src_valid),                                                  //          .valid
		.src_data           (id_router_012_src_data),                                                   //          .data
		.src_channel        (id_router_012_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                             //          .endofpacket
	);

	system_0_id_router_004 id_router_013 (
		.sink_ready         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                              //       src.ready
		.src_valid          (id_router_013_src_valid),                                              //          .valid
		.src_data           (id_router_013_src_data),                                               //          .data
		.src_channel        (id_router_013_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                         //          .endofpacket
	);

	system_0_id_router_004 id_router_014 (
		.sink_ready         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                              //       src.ready
		.src_valid          (id_router_014_src_valid),                                              //          .valid
		.src_data           (id_router_014_src_data),                                               //          .data
		.src_channel        (id_router_014_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                         //          .endofpacket
	);

	system_0_id_router_004 id_router_015 (
		.sink_ready         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                              //       src.ready
		.src_valid          (id_router_015_src_valid),                                              //          .valid
		.src_data           (id_router_015_src_data),                                               //          .data
		.src_channel        (id_router_015_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                         //          .endofpacket
	);

	system_0_id_router_004 id_router_016 (
		.sink_ready         (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (isp1362_dc_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                               //       src.ready
		.src_valid          (id_router_016_src_valid),                                               //          .valid
		.src_data           (id_router_016_src_data),                                                //          .data
		.src_channel        (id_router_016_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_004 id_router_017 (
		.sink_ready         (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (isp1362_hc_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                               //       src.ready
		.src_valid          (id_router_017_src_valid),                                               //          .valid
		.src_data           (id_router_017_src_data),                                                //          .data
		.src_channel        (id_router_017_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_004 id_router_018 (
		.sink_ready         (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                         //       src.ready
		.src_valid          (id_router_018_src_valid),                                                         //          .valid
		.src_data           (id_router_018_src_data),                                                          //          .data
		.src_channel        (id_router_018_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                    //          .endofpacket
	);

	system_0_id_router_004 id_router_019 (
		.sink_ready         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                           //       src.ready
		.src_valid          (id_router_019_src_valid),                                                           //          .valid
		.src_data           (id_router_019_src_data),                                                            //          .data
		.src_channel        (id_router_019_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                                      //          .endofpacket
	);

	system_0_id_router_004 id_router_020 (
		.sink_ready         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seg7_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                      //       src.ready
		.src_valid          (id_router_020_src_valid),                                                      //          .valid
		.src_data           (id_router_020_src_data),                                                       //          .data
		.src_channel        (id_router_020_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                                 //          .endofpacket
	);

	system_0_id_router_021 id_router_021 (
		.sink_ready         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                          //       src.ready
		.src_valid          (id_router_021_src_valid),                                                          //          .valid
		.src_data           (id_router_021_src_data),                                                           //          .data
		.src_channel        (id_router_021_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                                     //          .endofpacket
	);

	system_0_id_router_004 id_router_022 (
		.sink_ready         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                               //       src.ready
		.src_valid          (id_router_022_src_valid),                                               //          .valid
		.src_data           (id_router_022_src_data),                                                //          .data
		.src_channel        (id_router_022_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_004 id_router_023 (
		.sink_ready         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                               //       src.ready
		.src_valid          (id_router_023_src_valid),                                               //          .valid
		.src_data           (id_router_023_src_data),                                                //          .data
		.src_channel        (id_router_023_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_004 id_router_024 (
		.sink_ready         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_wp_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                               //       src.ready
		.src_valid          (id_router_024_src_valid),                                               //          .valid
		.src_data           (id_router_024_src_data),                                                //          .data
		.src_channel        (id_router_024_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_004 id_router_025 (
		.sink_ready         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_audio_clk_in_clk),                                                          //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                       //       src.ready
		.src_valid          (id_router_025_src_valid),                                                       //          .valid
		.src_data           (id_router_025_src_data),                                                        //          .data
		.src_channel        (id_router_025_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                                  //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (62),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (26),
		.VALID_WIDTH               (26),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (45),
		.PKT_BYTE_CNT_H            (41),
		.PKT_BYTE_CNT_L            (39),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (44),
		.PKT_BURSTWRAP_L           (42),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.ST_DATA_W                 (57),
		.ST_CHANNEL_W              (26),
		.OUT_BYTE_CNT_H            (39),
		.OUT_BURSTWRAP_H           (44),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),         //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),          //          .data
		.sink0_channel         (width_adapter_002_src_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),         //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (54),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (26),
		.OUT_BYTE_CNT_H            (49),
		.OUT_BURSTWRAP_H           (53),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (clk),                                     //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),                 //     sink0.valid
		.sink0_data            (width_adapter_src_data),                  //          .data
		.sink0_channel         (width_adapter_src_channel),               //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),         //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),           //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),                 //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (54),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (26),
		.OUT_BYTE_CNT_H            (49),
		.OUT_BURSTWRAP_H           (53),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_002 (
		.clk                   (clk),                                     //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_n),                            // reset_in0.reset
		.reset_in1  (~reset_n),                            // reset_in1.reset
		.reset_in2  (cpu_0_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (clk),                                 //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (~reset_n),                           // reset_in1.reset
		.clk        (clk),                                //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (~reset_n),                           // reset_in1.reset
		.clk        (clk_audio_clk_in_clk),               //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("none"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_n), // reset_in0.reset
		.reset_in1  (~reset_n), // reset_in1.reset
		.clk        (),         //       clk.clk
		.reset_out  (),         // reset_out.reset
		.reset_in2  (1'b0),     // (terminated)
		.reset_in3  (1'b0),     // (terminated)
		.reset_in4  (1'b0),     // (terminated)
		.reset_in5  (1'b0),     // (terminated)
		.reset_in6  (1'b0),     // (terminated)
		.reset_in7  (1'b0),     // (terminated)
		.reset_in8  (1'b0),     // (terminated)
		.reset_in9  (1'b0),     // (terminated)
		.reset_in10 (1'b0),     // (terminated)
		.reset_in11 (1'b0),     // (terminated)
		.reset_in12 (1'b0),     // (terminated)
		.reset_in13 (1'b0),     // (terminated)
		.reset_in14 (1'b0),     // (terminated)
		.reset_in15 (1'b0)      // (terminated)
	);

	system_0_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk),                               //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)    //           .endofpacket
	);

	system_0_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk),                                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_001_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_001_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_001_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_001_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_001_src22_endofpacket),   //          .endofpacket
		.src23_ready         (cmd_xbar_demux_001_src23_ready),         //     src23.ready
		.src23_valid         (cmd_xbar_demux_001_src23_valid),         //          .valid
		.src23_data          (cmd_xbar_demux_001_src23_data),          //          .data
		.src23_channel       (cmd_xbar_demux_001_src23_channel),       //          .channel
		.src23_startofpacket (cmd_xbar_demux_001_src23_startofpacket), //          .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_001_src23_endofpacket),   //          .endofpacket
		.src24_ready         (cmd_xbar_demux_001_src24_ready),         //     src24.ready
		.src24_valid         (cmd_xbar_demux_001_src24_valid),         //          .valid
		.src24_data          (cmd_xbar_demux_001_src24_data),          //          .data
		.src24_channel       (cmd_xbar_demux_001_src24_channel),       //          .channel
		.src24_startofpacket (cmd_xbar_demux_001_src24_startofpacket), //          .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_001_src24_endofpacket),   //          .endofpacket
		.src25_ready         (cmd_xbar_demux_001_src25_ready),         //     src25.ready
		.src25_valid         (cmd_xbar_demux_001_src25_valid),         //          .valid
		.src25_data          (cmd_xbar_demux_001_src25_data),          //          .data
		.src25_channel       (cmd_xbar_demux_001_src25_channel),       //          .channel
		.src25_startofpacket (cmd_xbar_demux_001_src25_startofpacket), //          .startofpacket
		.src25_endofpacket   (cmd_xbar_demux_001_src25_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk),                                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk),                                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk),                                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk),                                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_005 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_006 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_007 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_008 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_009 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_010 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_011 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_012 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_013 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_014 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_015 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_016 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_017 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_018 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_019 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_020 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_021 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_005_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_005_src_channel),         //          .channel
		.sink_data          (width_adapter_005_src_data),            //          .data
		.sink_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_005_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_022 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_023 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_024 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_004 rsp_xbar_demux_025 (
		.clk                (clk_audio_clk_in_clk),                  //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk),                                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk),                                   //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_022_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_023_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_024_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink25_ready         (crosser_001_out_ready),                 //    sink25.ready
		.sink25_valid         (crosser_001_out_valid),                 //          .valid
		.sink25_channel       (crosser_001_out_channel),               //          .channel
		.sink25_data          (crosser_001_out_data),                  //          .data
		.sink25_startofpacket (crosser_001_out_startofpacket),         //          .startofpacket
		.sink25_endofpacket   (crosser_001_out_endofpacket)            //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (68),
		.IN_PKT_BYTE_CNT_L             (66),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (69),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (50),
		.OUT_PKT_BYTE_CNT_L            (48),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (26),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk               (clk),                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid          (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel        (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data           (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket   (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data          (width_adapter_src_data),             //          .data
		.out_channel       (width_adapter_src_channel),          //          .channel
		.out_valid         (width_adapter_src_valid),            //          .valid
		.out_ready         (width_adapter_src_ready),            //          .ready
		.out_startofpacket (width_adapter_src_startofpacket)     //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (50),
		.IN_PKT_BYTE_CNT_L             (48),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (53),
		.IN_PKT_BURSTWRAP_L            (51),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (68),
		.OUT_PKT_BYTE_CNT_L            (66),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (26),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk               (clk),                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid          (id_router_001_src_valid),             //      sink.valid
		.in_channel        (id_router_001_src_channel),           //          .channel
		.in_startofpacket  (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_001_src_ready),             //          .ready
		.in_data           (id_router_001_src_data),              //          .data
		.out_endofpacket   (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_001_src_data),          //          .data
		.out_channel       (width_adapter_001_src_channel),       //          .channel
		.out_valid         (width_adapter_001_src_valid),         //          .valid
		.out_ready         (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket (width_adapter_001_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (68),
		.IN_PKT_BYTE_CNT_L             (66),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (69),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (33),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (41),
		.OUT_PKT_BYTE_CNT_L            (39),
		.OUT_PKT_TRANS_COMPRESSED_READ (34),
		.OUT_ST_DATA_W                 (57),
		.ST_CHANNEL_W                  (26),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk               (clk),                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid          (cmd_xbar_mux_003_src_valid),          //      sink.valid
		.in_channel        (cmd_xbar_mux_003_src_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_mux_003_src_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_003_src_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_mux_003_src_ready),          //          .ready
		.in_data           (cmd_xbar_mux_003_src_data),           //          .data
		.out_endofpacket   (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_002_src_data),          //          .data
		.out_channel       (width_adapter_002_src_channel),       //          .channel
		.out_valid         (width_adapter_002_src_valid),         //          .valid
		.out_ready         (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket (width_adapter_002_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (33),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (41),
		.IN_PKT_BYTE_CNT_L             (39),
		.IN_PKT_TRANS_COMPRESSED_READ  (34),
		.IN_PKT_BURSTWRAP_H            (44),
		.IN_PKT_BURSTWRAP_L            (42),
		.IN_ST_DATA_W                  (57),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (68),
		.OUT_PKT_BYTE_CNT_L            (66),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (26),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk               (clk),                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid          (id_router_003_src_valid),             //      sink.valid
		.in_channel        (id_router_003_src_channel),           //          .channel
		.in_startofpacket  (id_router_003_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_003_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_003_src_ready),             //          .ready
		.in_data           (id_router_003_src_data),              //          .data
		.out_endofpacket   (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_003_src_data),          //          .data
		.out_channel       (width_adapter_003_src_channel),       //          .channel
		.out_valid         (width_adapter_003_src_valid),         //          .valid
		.out_ready         (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket (width_adapter_003_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (68),
		.IN_PKT_BYTE_CNT_L             (66),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (69),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (50),
		.OUT_PKT_BYTE_CNT_L            (48),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (26),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_004 (
		.clk               (clk),                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_001_src21_valid),         //      sink.valid
		.in_channel        (cmd_xbar_demux_001_src21_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src21_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_demux_001_src21_ready),         //          .ready
		.in_data           (cmd_xbar_demux_001_src21_data),          //          .data
		.out_endofpacket   (width_adapter_004_src_endofpacket),      //       src.endofpacket
		.out_data          (width_adapter_004_src_data),             //          .data
		.out_channel       (width_adapter_004_src_channel),          //          .channel
		.out_valid         (width_adapter_004_src_valid),            //          .valid
		.out_ready         (width_adapter_004_src_ready),            //          .ready
		.out_startofpacket (width_adapter_004_src_startofpacket)     //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (50),
		.IN_PKT_BYTE_CNT_L             (48),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (53),
		.IN_PKT_BURSTWRAP_L            (51),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (68),
		.OUT_PKT_BYTE_CNT_L            (66),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (26),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_005 (
		.clk               (clk),                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid          (id_router_021_src_valid),             //      sink.valid
		.in_channel        (id_router_021_src_channel),           //          .channel
		.in_startofpacket  (id_router_021_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_021_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_021_src_ready),             //          .ready
		.in_data           (id_router_021_src_data),              //          .data
		.out_endofpacket   (width_adapter_005_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_005_src_data),          //          .data
		.out_channel       (width_adapter_005_src_channel),       //          .channel
		.out_valid         (width_adapter_005_src_valid),         //          .valid
		.out_ready         (width_adapter_005_src_ready),         //          .ready
		.out_startofpacket (width_adapter_005_src_startofpacket)  //          .startofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (84),
		.BITS_PER_SYMBOL     (84),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (26),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk),                                    //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (clk_audio_clk_in_clk),                   //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src25_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src25_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src25_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src25_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src25_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src25_data),          //              .data
		.out_ready         (crosser_out_ready),                      //           out.ready
		.out_valid         (crosser_out_valid),                      //              .valid
		.out_startofpacket (crosser_out_startofpacket),              //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),                //              .endofpacket
		.out_channel       (crosser_out_channel),                    //              .channel
		.out_data          (crosser_out_data),                       //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (84),
		.BITS_PER_SYMBOL     (84),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (26),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_audio_clk_in_clk),                  //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk),                                   //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_025_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_025_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_025_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_025_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_025_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_025_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	system_0_irq_mapper irq_mapper (
		.clk           (clk),                            //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (~irq_mapper_receiver7_irq),      // receiver7.irq
		.receiver8_irq (~irq_mapper_receiver8_irq),      // receiver8.irq
		.sender_irq    (cpu_0_d_irq_irq)                 //    sender.irq
	);

endmodule
