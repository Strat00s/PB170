library verilog;
use verilog.vl_types.all;
entity knight_rider_vlg_sample_tst is
    port(
        CLOCK_50        : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end knight_rider_vlg_sample_tst;
