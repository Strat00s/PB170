library verilog;
use verilog.vl_types.all;
entity knight_rider_vlg_vec_tst is
end knight_rider_vlg_vec_tst;
