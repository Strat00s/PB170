library verilog;
use verilog.vl_types.all;
entity PWM is
    port(
        clk             : in     vl_logic;
        \out\           : out    vl_logic
    );
end PWM;
